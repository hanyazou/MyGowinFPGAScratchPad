module sseg_decoder(
   input wire logic [3:0] num,
   output reg [6:0] y
   );

   /*
    *           A
    *         -----
    *      F/  G  /B
    *       -----
    *    E/     /C
    *     -----
    *       D
    */

   always_comb begin
      case (num)       // GFE DCBA
        4'b0000  : y = 7'b100_0000;  // 0
        4'b0001  : y = 7'b111_1001;  // 1
        4'b0010  : y = 7'b010_0100;  // 2
        4'b0011  : y = 7'b011_0000;  // 3
        4'b0100  : y = 7'b001_1001;  // 4
        4'b0101  : y = 7'b001_0010;  // 5
        4'b0110  : y = 7'b000_0010;  // 6
        4'b0111  : y = 7'b101_1000;  // 7
        4'b1000  : y = 7'b000_0000;  // 8
        4'b1001  : y = 7'b001_0000;  // 9
        4'b1010  : y = 7'b000_1000;  // A
        4'b1011  : y = 7'b000_0011;  // b
        4'b1100  : y = 7'b100_0110;  // C
        4'b1101  : y = 7'b010_0001;  // d
        4'b1110  : y = 7'b000_0110;  // E
        4'b1111  : y = 7'b000_1110;  // F
      endcase
   end

endmodule  // sseg_decoder
