   `include "h80cpu.svh"
   `include "h80cpu_instmacros.svh"
   initial begin
      mem0[16'h0000]=16'h0160;
      mem1[16'h0000]=16'h0100;
      mem0[16'h0001]=16'h01e0;
      mem1[16'h0001]=16'hffff;
      mem0[16'h0002]=16'hffff;
      mem1[16'h0002]=16'hffff;
      mem0[16'h0003]=16'hffff;
      mem1[16'h0003]=16'hffff;
      mem0[16'h0004]=16'h0160;
      mem1[16'h0004]=16'h0ab8;
      mem0[16'h0005]=16'h01e0;
      mem1[16'h0005]=16'hffff;
      mem0[16'h0006]=16'h0160;
      mem1[16'h0006]=16'h0ad4;
      mem0[16'h0007]=16'h01e0;
      mem1[16'h0007]=16'hffff;
      mem0[16'h0008]=16'hffff;
      mem1[16'h0008]=16'hffff;
      mem0[16'h0009]=16'hffff;
      mem1[16'h0009]=16'hffff;
      mem0[16'h000a]=16'hffff;
      mem1[16'h000a]=16'hffff;
      mem0[16'h000b]=16'hffff;
      mem1[16'h000b]=16'hffff;
      mem0[16'h000c]=16'h0160;
      mem1[16'h000c]=16'h0a32;
      mem0[16'h000d]=16'h01e0;
      mem1[16'h000d]=16'hffff;
      mem0[16'h000e]=16'h0160;
      mem1[16'h000e]=16'h0a34;
      mem0[16'h000f]=16'h01e0;
      mem1[16'h000f]=16'hffff;
      mem0[16'h0010]=16'hffff;
      mem1[16'h0010]=16'hffff;
      mem0[16'h0011]=16'hffff;
      mem1[16'h0011]=16'hffff;
      mem0[16'h0012]=16'hffff;
      mem1[16'h0012]=16'hffff;
      mem0[16'h0013]=16'hffff;
      mem1[16'h0013]=16'hffff;
      mem0[16'h0014]=16'hffff;
      mem1[16'h0014]=16'hffff;
      mem0[16'h0015]=16'hffff;
      mem1[16'h0015]=16'hffff;
      mem0[16'h0016]=16'hffff;
      mem1[16'h0016]=16'hffff;
      mem0[16'h0017]=16'hffff;
      mem1[16'h0017]=16'hffff;
      mem0[16'h0018]=16'hffff;
      mem1[16'h0018]=16'hffff;
      mem0[16'h0019]=16'hffff;
      mem1[16'h0019]=16'hffff;
      mem0[16'h001a]=16'hffff;
      mem1[16'h001a]=16'hffff;
      mem0[16'h001b]=16'hffff;
      mem1[16'h001b]=16'hffff;
      mem0[16'h001c]=16'hffff;
      mem1[16'h001c]=16'hffff;
      mem0[16'h001d]=16'hffff;
      mem1[16'h001d]=16'hffff;
      mem0[16'h001e]=16'hffff;
      mem1[16'h001e]=16'hffff;
      mem0[16'h001f]=16'hffff;
      mem1[16'h001f]=16'hffff;
      mem0[16'h0020]=16'h0160;
      mem1[16'h0020]=16'h0100;
      mem0[16'h0021]=16'h01e0;
      mem1[16'h0021]=16'hffff;
      mem0[16'h0022]=16'h0160;
      mem1[16'h0022]=16'h01fc;
      mem0[16'h0023]=16'h01e0;
      mem1[16'h0023]=16'hffff;
      mem0[16'h0024]=16'h0160;
      mem1[16'h0024]=16'h0ad4;
      mem0[16'h0025]=16'h01e0;
      mem1[16'h0025]=16'hffff;
      mem0[16'h0026]=16'h0160;
      mem1[16'h0026]=16'h087c;
      mem0[16'h0027]=16'h01e0;
      mem1[16'h0027]=16'hffff;
      mem0[16'h0028]=16'h0160;
      mem1[16'h0028]=16'h0ab8;
      mem0[16'h0029]=16'h01e0;
      mem1[16'h0029]=16'hffff;
      mem0[16'h002a]=16'h0160;
      mem1[16'h002a]=16'h0aca;
      mem0[16'h002b]=16'h01e0;
      mem1[16'h002b]=16'hffff;
      mem0[16'h002c]=16'hffff;
      mem1[16'h002c]=16'hffff;
      mem0[16'h002d]=16'hffff;
      mem1[16'h002d]=16'hffff;
      mem0[16'h002e]=16'hffff;
      mem1[16'h002e]=16'hffff;
      mem0[16'h002f]=16'hffff;
      mem1[16'h002f]=16'hffff;
      mem0[16'h0030]=16'hffff;
      mem1[16'h0030]=16'hffff;
      mem0[16'h0031]=16'hffff;
      mem1[16'h0031]=16'hffff;
      mem0[16'h0032]=16'hffff;
      mem1[16'h0032]=16'hffff;
      mem0[16'h0033]=16'hffff;
      mem1[16'h0033]=16'hffff;
      mem0[16'h0034]=16'hffff;
      mem1[16'h0034]=16'hffff;
      mem0[16'h0035]=16'hffff;
      mem1[16'h0035]=16'hffff;
      mem0[16'h0036]=16'hffff;
      mem1[16'h0036]=16'hffff;
      mem0[16'h0037]=16'hffff;
      mem1[16'h0037]=16'hffff;
      mem0[16'h0038]=16'hffff;
      mem1[16'h0038]=16'hffff;
      mem0[16'h0039]=16'hffff;
      mem1[16'h0039]=16'hffff;
      mem0[16'h003a]=16'hffff;
      mem1[16'h003a]=16'hffff;
      mem0[16'h003b]=16'hffff;
      mem1[16'h003b]=16'hffff;
      mem0[16'h003c]=16'hffff;
      mem1[16'h003c]=16'hffff;
      mem0[16'h003d]=16'hffff;
      mem1[16'h003d]=16'hffff;
      mem0[16'h003e]=16'hffff;
      mem1[16'h003e]=16'hffff;
      mem0[16'h003f]=16'hffff;
      mem1[16'h003f]=16'hffff;
      mem0[16'h0040]=16'h0166;
      mem1[16'h0040]=16'h0ff0;
      mem0[16'h0041]=16'h3f26;
      mem1[16'h0041]=16'h0169;
      mem0[16'h0042]=16'h1000;
      mem1[16'h0042]=16'h016a;
      mem0[16'h0043]=16'h1001;
      mem1[16'h0043]=16'he666;
      mem0[16'h0044]=16'he777;
      mem1[16'h0044]=16'h3a6a;
      mem0[16'h0045]=16'h3c67;
      mem1[16'h0045]=16'h0146;
      mem0[16'h0046]=16'h10ff;
      mem1[16'h0046]=16'hc660;
      mem0[16'h0047]=16'h386a;
      mem1[16'h0047]=16'h3a4a;
      mem0[16'h0048]=16'hf664;
      mem1[16'h0048]=16'h0170;
      mem0[16'h0049]=16'h001a;
      mem1[16'h0049]=16'h0380;
      mem0[16'h004a]=16'h3a69;
      mem1[16'h004a]=16'hf664;
      mem0[16'h004b]=16'h0170;
      mem1[16'h004b]=16'h001c;
      mem0[16'h004c]=16'h0380;
      mem1[16'h004c]=16'h387a;
      mem0[16'h004d]=16'h3a69;
      mem1[16'h004d]=16'h3a4a;
      mem0[16'h004e]=16'hf664;
      mem1[16'h004e]=16'h0170;
      mem0[16'h004f]=16'h000e;
      mem1[16'h004f]=16'h0380;
      mem0[16'h0050]=16'h0160;
      mem1[16'h0050]=16'h0f20;
      mem0[16'h0051]=16'h34a0;
      mem1[16'h0051]=16'h0170;
      mem0[16'h0052]=16'h001a;
      mem1[16'h0052]=16'h01f0;
      mem0[16'h0053]=16'h387a;
      mem1[16'h0053]=16'h08a1;
      mem0[16'h0054]=16'h00f0;
      mem1[16'h0054]=16'h0000;
      mem0[16'h0055]=16'h0001;
      mem1[16'h0055]=16'hfaa0;
      mem0[16'h0056]=16'h0170;
      mem1[16'h0056]=16'hffb6;
      mem0[16'h0057]=16'h0380;
      mem1[16'h0057]=16'h0160;
      mem0[16'h0058]=16'h0f20;
      mem1[16'h0058]=16'h34a0;
      mem0[16'h0059]=16'he666;
      mem1[16'h0059]=16'h0160;
      mem0[16'h005a]=16'h0f1c;
      mem1[16'h005a]=16'h3860;
      mem0[16'h005b]=16'h0168;
      mem1[16'h005b]=16'h0aa1;
      mem0[16'h005c]=16'he999;
      mem1[16'h005c]=16'h0160;
      mem0[16'h005d]=16'h0178;
      mem1[16'h005d]=16'h01e0;
      mem0[16'h005e]=16'h0160;
      mem1[16'h005e]=16'h0f1c;
      mem0[16'h005f]=16'h3890;
      mem1[16'h005f]=16'h0160;
      mem0[16'h0060]=16'h0f00;
      mem1[16'h0060]=16'h3480;
      mem0[16'h0061]=16'h0160;
      mem1[16'h0061]=16'h0ab6;
      mem0[16'h0062]=16'h01c0;
      mem1[16'h0062]=16'h0166;
      mem0[16'h0063]=16'h1000;
      mem1[16'h0063]=16'h0160;
      mem0[16'h0064]=16'h0f10;
      mem1[16'h0064]=16'h3460;
      mem0[16'h0065]=16'h0160;
      mem1[16'h0065]=16'h0f18;
      mem0[16'h0066]=16'h3460;
      mem1[16'h0066]=16'h0160;
      mem0[16'h0067]=16'h0f16;
      mem1[16'h0067]=16'h3460;
      mem0[16'h0068]=16'h1649;
      mem1[16'h0068]=16'h0160;
      mem0[16'h0069]=16'h0f1a;
      mem1[16'h0069]=16'h3860;
      mem0[16'h006a]=16'he666;
      mem1[16'h006a]=16'h0160;
      mem0[16'h006b]=16'h0f1e;
      mem1[16'h006b]=16'h3860;
      mem0[16'h006c]=16'h1864;
      mem1[16'h006c]=16'he222;
      mem0[16'h006d]=16'h0160;
      mem1[16'h006d]=16'h0ad4;
      mem0[16'h006e]=16'h01c0;
      mem1[16'h006e]=16'h0170;
      mem0[16'h006f]=16'hfff4;
      mem1[16'h006f]=16'h0a80;
      mem0[16'h0070]=16'h0164;
      mem1[16'h0070]=16'h0a36;
      mem0[16'h0071]=16'h0160;
      mem1[16'h0071]=16'h087c;
      mem0[16'h0072]=16'h01c0;
      mem1[16'h0072]=16'h0160;
      mem0[16'h0073]=16'h0f00;
      mem1[16'h0073]=16'h3640;
      mem0[16'h0074]=16'h0160;
      mem1[16'h0074]=16'h087c;
      mem0[16'h0075]=16'h01c0;
      mem1[16'h0075]=16'h0164;
      mem0[16'h0076]=16'h1000;
      mem1[16'h0076]=16'h0160;
      mem0[16'h0077]=16'h0890;
      mem1[16'h0077]=16'h01c0;
      mem0[16'h0078]=16'h122d;
      mem1[16'h0078]=16'h0160;
      mem0[16'h0079]=16'h0ad4;
      mem1[16'h0079]=16'h01c0;
      mem0[16'h007a]=16'h0160;
      mem1[16'h007a]=16'h0f20;
      mem0[16'h007b]=16'h3640;
      mem1[16'h007b]=16'h0941;
      mem0[16'h007c]=16'h0160;
      mem1[16'h007c]=16'h0890;
      mem0[16'h007d]=16'h01c0;
      mem1[16'h007d]=16'h0160;
      mem0[16'h007e]=16'h0910;
      mem1[16'h007e]=16'h01c0;
      mem0[16'h007f]=16'h0164;
      mem1[16'h007f]=16'h0a50;
      mem0[16'h0080]=16'h0160;
      mem1[16'h0080]=16'h087c;
      mem0[16'h0081]=16'h01c0;
      mem1[16'h0081]=16'h0160;
      mem0[16'h0082]=16'h0920;
      mem1[16'h0082]=16'h01c0;
      mem0[16'h0083]=16'h0164;
      mem1[16'h0083]=16'h0f00;
      mem0[16'h0084]=16'h0160;
      mem1[16'h0084]=16'h09c2;
      mem0[16'h0085]=16'h01c0;
      mem1[16'h0085]=16'h0160;
      mem0[16'h0086]=16'h09d4;
      mem1[16'h0086]=16'h01c0;
      mem0[16'h0087]=16'hd222;
      mem1[16'h0087]=16'h0170;
      mem0[16'h0088]=16'hffda;
      mem1[16'h0088]=16'h03c0;
      mem0[16'h0089]=16'h1044;
      mem1[16'h0089]=16'hf220;
      mem0[16'h008a]=16'h0170;
      mem1[16'h008a]=16'h003a;
      mem0[16'h008b]=16'h03c0;
      mem1[16'h008b]=16'h1047;
      mem0[16'h008c]=16'hf220;
      mem1[16'h008c]=16'h0160;
      mem0[16'h008d]=16'h0444;
      mem1[16'h008d]=16'h0340;
      mem0[16'h008e]=16'h1053;
      mem1[16'h008e]=16'hf220;
      mem0[16'h008f]=16'h0160;
      mem1[16'h008f]=16'h0476;
      mem0[16'h0090]=16'h0340;
      mem1[16'h0090]=16'h104c;
      mem0[16'h0091]=16'hf220;
      mem1[16'h0091]=16'h0160;
      mem0[16'h0092]=16'h0544;
      mem1[16'h0092]=16'h0340;
      mem0[16'h0093]=16'h1050;
      mem1[16'h0093]=16'hf220;
      mem0[16'h0094]=16'h0160;
      mem1[16'h0094]=16'h06ea;
      mem0[16'h0095]=16'h0340;
      mem1[16'h0095]=16'h0164;
      mem0[16'h0096]=16'h0a6d;
      mem1[16'h0096]=16'h0160;
      mem0[16'h0097]=16'h087c;
      mem1[16'h0097]=16'h01c0;
      mem0[16'h0098]=16'h0170;
      mem1[16'h0098]=16'hff98;
      mem0[16'h0099]=16'h01f0;
      mem1[16'h0099]=16'h0841;
      mem0[16'h009a]=16'h0160;
      mem1[16'h009a]=16'h09c2;
      mem0[16'h009b]=16'h01c0;
      mem1[16'h009b]=16'h0160;
      mem0[16'h009c]=16'h09e6;
      mem1[16'h009c]=16'h01c0;
      mem0[16'h009d]=16'hd333;
      mem1[16'h009d]=16'h0170;
      mem0[16'h009e]=16'h0026;
      mem1[16'h009e]=16'h0380;
      mem0[16'h009f]=16'h0160;
      mem1[16'h009f]=16'h09c2;
      mem0[16'h00a0]=16'h01c0;
      mem1[16'h00a0]=16'hd222;
      mem0[16'h00a1]=16'h0170;
      mem1[16'h00a1]=16'hffce;
      mem0[16'h00a2]=16'h0380;
      mem1[16'h00a2]=16'h0160;
      mem0[16'h00a3]=16'h0f10;
      mem1[16'h00a3]=16'h3660;
      mem0[16'h00a4]=16'h1080;
      mem1[16'h00a4]=16'h8660;
      mem0[16'h00a5]=16'h0160;
      mem1[16'h00a5]=16'h0f12;
      mem0[16'h00a6]=16'h3460;
      mem1[16'h00a6]=16'h0170;
      mem0[16'h00a7]=16'h005c;
      mem1[16'h00a7]=16'h01f0;
      mem0[16'h00a8]=16'h0160;
      mem1[16'h00a8]=16'h0f10;
      mem0[16'h00a9]=16'h3450;
      mem1[16'h00a9]=16'h0160;
      mem0[16'h00aa]=16'h09c2;
      mem1[16'h00aa]=16'h01c0;
      mem0[16'h00ab]=16'h102c;
      mem1[16'h00ab]=16'hf220;
      mem0[16'h00ac]=16'h0170;
      mem1[16'h00ac]=16'h001a;
      mem0[16'h00ad]=16'h03c0;
      mem1[16'h00ad]=16'hd222;
      mem0[16'h00ae]=16'h0170;
      mem1[16'h00ae]=16'hff9a;
      mem0[16'h00af]=16'h0380;
      mem1[16'h00af]=16'h1080;
      mem0[16'h00b0]=16'h8550;
      mem1[16'h00b0]=16'h0160;
      mem0[16'h00b1]=16'h0f12;
      mem1[16'h00b1]=16'h3450;
      mem0[16'h00b2]=16'h0170;
      mem1[16'h00b2]=16'h002e;
      mem0[16'h00b3]=16'h01f0;
      mem1[16'h00b3]=16'h0841;
      mem0[16'h00b4]=16'h0160;
      mem1[16'h00b4]=16'h09c2;
      mem0[16'h00b5]=16'h01c0;
      mem1[16'h00b5]=16'h0160;
      mem0[16'h00b6]=16'h09e6;
      mem1[16'h00b6]=16'h01c0;
      mem0[16'h00b7]=16'h0160;
      mem1[16'h00b7]=16'h09c2;
      mem0[16'h00b8]=16'h01c0;
      mem1[16'h00b8]=16'hd333;
      mem0[16'h00b9]=16'h0170;
      mem1[16'h00b9]=16'hff6e;
      mem0[16'h00ba]=16'h03c0;
      mem1[16'h00ba]=16'hd222;
      mem0[16'h00bb]=16'h0160;
      mem1[16'h00bb]=16'h0256;
      mem0[16'h00bc]=16'h0300;
      mem1[16'h00bc]=16'h0851;
      mem0[16'h00bd]=16'h0160;
      mem1[16'h00bd]=16'h0f12;
      mem0[16'h00be]=16'h3450;
      mem1[16'h00be]=16'he444;
      mem0[16'h00bf]=16'h0160;
      mem1[16'h00bf]=16'h0f10;
      mem0[16'h00c0]=16'h3640;
      mem1[16'h00c0]=16'h0160;
      mem0[16'h00c1]=16'hfff0;
      mem1[16'h00c1]=16'hc440;
      mem0[16'h00c2]=16'he666;
      mem1[16'h00c2]=16'h0160;
      mem0[16'h00c3]=16'h0f14;
      mem1[16'h00c3]=16'h3860;
      mem0[16'h00c4]=16'h0104;
      mem1[16'h00c4]=16'h0160;
      mem0[16'h00c5]=16'h035e;
      mem1[16'h00c5]=16'h01c0;
      mem0[16'h00c6]=16'h0114;
      mem1[16'h00c6]=16'h1010;
      mem0[16'h00c7]=16'h8440;
      mem1[16'h00c7]=16'h0160;
      mem0[16'h00c8]=16'h0aca;
      mem1[16'h00c8]=16'h01c0;
      mem0[16'h00c9]=16'h0170;
      mem1[16'h00c9]=16'h0024;
      mem0[16'h00ca]=16'h0380;
      mem1[16'h00ca]=16'h0160;
      mem0[16'h00cb]=16'h0f14;
      mem1[16'h00cb]=16'h3a20;
      mem0[16'h00cc]=16'h1002;
      mem1[16'h00cc]=16'hf220;
      mem0[16'h00cd]=16'h0170;
      mem1[16'h00cd]=16'hffd8;
      mem0[16'h00ce]=16'h03d0;
      mem1[16'h00ce]=16'h0160;
      mem0[16'h00cf]=16'h0f12;
      mem1[16'h00cf]=16'h3640;
      mem0[16'h00d0]=16'h0160;
      mem1[16'h00d0]=16'h0f10;
      mem0[16'h00d1]=16'h3440;
      mem1[16'h00d1]=16'h0160;
      mem0[16'h00d2]=16'h01fc;
      mem1[16'h00d2]=16'h01e0;
      mem0[16'h00d3]=16'h0160;
      mem1[16'h00d3]=16'h0f10;
      mem0[16'h00d4]=16'h3440;
      mem1[16'h00d4]=16'h0160;
      mem0[16'h00d5]=16'h0ab8;
      mem1[16'h00d5]=16'h01c0;
      mem0[16'h00d6]=16'h0160;
      mem1[16'h00d6]=16'h01fc;
      mem0[16'h00d7]=16'h01e0;
      mem1[16'h00d7]=16'h0160;
      mem0[16'h00d8]=16'h0890;
      mem1[16'h00d8]=16'h01c0;
      mem0[16'h00d9]=16'h0104;
      mem1[16'h00d9]=16'h0164;
      mem0[16'h00da]=16'h0a75;
      mem1[16'h00da]=16'h0160;
      mem0[16'h00db]=16'h087c;
      mem1[16'h00db]=16'h01c0;
      mem0[16'h00dc]=16'h0114;
      mem1[16'h00dc]=16'h0168;
      mem0[16'h00dd]=16'h0f00;
      mem1[16'h00dd]=16'h1910;
      mem0[16'h00de]=16'h0160;
      mem1[16'h00de]=16'h03cc;
      mem0[16'h00df]=16'h01c0;
      mem1[16'h00df]=16'h0170;
      mem0[16'h00e0]=16'hfff6;
      mem1[16'h00e0]=16'h0a90;
      mem0[16'h00e1]=16'h0164;
      mem1[16'h00e1]=16'h0a78;
      mem0[16'h00e2]=16'h0160;
      mem1[16'h00e2]=16'h087c;
      mem0[16'h00e3]=16'h01c0;
      mem1[16'h00e3]=16'h0164;
      mem0[16'h00e4]=16'h0f00;
      mem1[16'h00e4]=16'h1910;
      mem0[16'h00e5]=16'h3a24;
      mem1[16'h00e5]=16'h0841;
      mem0[16'h00e6]=16'h1020;
      mem1[16'h00e6]=16'hf220;
      mem0[16'h00e7]=16'h0170;
      mem1[16'h00e7]=16'h0018;
      mem0[16'h00e8]=16'h03d0;
      mem1[16'h00e8]=16'h107f;
      mem0[16'h00e9]=16'hf220;
      mem1[16'h00e9]=16'h0170;
      mem0[16'h00ea]=16'h000e;
      mem1[16'h00ea]=16'h0390;
      mem0[16'h00eb]=16'h0160;
      mem1[16'h00eb]=16'h0ad4;
      mem0[16'h00ec]=16'h01c0;
      mem1[16'h00ec]=16'h0170;
      mem0[16'h00ed]=16'h000a;
      mem1[16'h00ed]=16'h01f0;
      mem0[16'h00ee]=16'h122e;
      mem1[16'h00ee]=16'h0160;
      mem0[16'h00ef]=16'h0ad4;
      mem1[16'h00ef]=16'h01c0;
      mem0[16'h00f0]=16'h0170;
      mem1[16'h00f0]=16'hffd0;
      mem0[16'h00f1]=16'h0a90;
      mem1[16'h00f1]=16'h0160;
      mem0[16'h00f2]=16'h0910;
      mem1[16'h00f2]=16'h01e0;
      mem0[16'h00f3]=16'h1220;
      mem1[16'h00f3]=16'h0160;
      mem0[16'h00f4]=16'h0ad4;
      mem1[16'h00f4]=16'h01c0;
      mem0[16'h00f5]=16'he666;
      mem1[16'h00f5]=16'h0160;
      mem0[16'h00f6]=16'h0f14;
      mem1[16'h00f6]=16'h3a60;
      mem0[16'h00f7]=16'hd666;
      mem1[16'h00f7]=16'h0170;
      mem0[16'h00f8]=16'h0030;
      mem1[16'h00f8]=16'h0380;
      mem0[16'h00f9]=16'he666;
      mem1[16'h00f9]=16'h0160;
      mem0[16'h00fa]=16'h0f10;
      mem1[16'h00fa]=16'h3660;
      mem0[16'h00fb]=16'hf664;
      mem1[16'h00fb]=16'h0170;
      mem0[16'h00fc]=16'h0018;
      mem1[16'h00fc]=16'h03c0;
      mem0[16'h00fd]=16'h1220;
      mem1[16'h00fd]=16'h0160;
      mem0[16'h00fe]=16'h0ad4;
      mem1[16'h00fe]=16'h01c0;
      mem0[16'h00ff]=16'h0160;
      mem1[16'h00ff]=16'h0ad4;
      mem0[16'h0100]=16'h01c0;
      mem1[16'h0100]=16'h3828;
      mem0[16'h0101]=16'h0841;
      mem1[16'h0101]=16'h0881;
      mem0[16'h0102]=16'h0002;
      mem1[16'h0102]=16'h1601;
      mem0[16'h0103]=16'h0160;
      mem1[16'h0103]=16'h0f14;
      mem0[16'h0104]=16'h3860;
      mem1[16'h0104]=16'h0160;
      mem0[16'h0105]=16'h0f14;
      mem1[16'h0105]=16'h3a60;
      mem0[16'h0106]=16'h1001;
      mem1[16'h0106]=16'hf660;
      mem0[16'h0107]=16'h0170;
      mem1[16'h0107]=16'hffd4;
      mem0[16'h0108]=16'h0380;
      mem1[16'h0108]=16'h3a24;
      mem0[16'h0109]=16'h3828;
      mem1[16'h0109]=16'h0160;
      mem0[16'h010a]=16'h089c;
      mem1[16'h010a]=16'h01c0;
      mem0[16'h010b]=16'h0841;
      mem1[16'h010b]=16'h0881;
      mem0[16'h010c]=16'h0160;
      mem1[16'h010c]=16'h0f12;
      mem0[16'h010d]=16'h3660;
      mem1[16'h010d]=16'hf446;
      mem0[16'h010e]=16'h0080;
      mem1[16'h010e]=16'h1602;
      mem0[16'h010f]=16'h0160;
      mem1[16'h010f]=16'h0f14;
      mem0[16'h0110]=16'h3860;
      mem1[16'h0110]=16'h0002;
      mem0[16'h0111]=16'h0841;
      mem1[16'h0111]=16'h0160;
      mem0[16'h0112]=16'h09c2;
      mem1[16'h0112]=16'h01c0;
      mem0[16'h0113]=16'h0160;
      mem1[16'h0113]=16'h09e6;
      mem0[16'h0114]=16'h01c0;
      mem1[16'h0114]=16'h0160;
      mem0[16'h0115]=16'h09c2;
      mem1[16'h0115]=16'h01c0;
      mem0[16'h0116]=16'hd222;
      mem1[16'h0116]=16'h0160;
      mem0[16'h0117]=16'h0256;
      mem1[16'h0117]=16'h0300;
      mem0[16'h0118]=16'hd333;
      mem1[16'h0118]=16'h0170;
      mem0[16'h0119]=16'h0008;
      mem1[16'h0119]=16'h03c0;
      mem0[16'h011a]=16'h0160;
      mem1[16'h011a]=16'h0f16;
      mem0[16'h011b]=16'h3450;
      mem1[16'h011b]=16'h0160;
      mem0[16'h011c]=16'h0f16;
      mem1[16'h011c]=16'h3660;
      mem0[16'h011d]=16'h01e6;
      mem1[16'h011d]=16'h0841;
      mem0[16'h011e]=16'h0160;
      mem1[16'h011e]=16'h09c2;
      mem0[16'h011f]=16'h01c0;
      mem1[16'h011f]=16'h0160;
      mem0[16'h0120]=16'h09e6;
      mem1[16'h0120]=16'h01c0;
      mem0[16'h0121]=16'h0160;
      mem1[16'h0121]=16'h09c2;
      mem0[16'h0122]=16'h01c0;
      mem1[16'h0122]=16'hd222;
      mem0[16'h0123]=16'h0160;
      mem1[16'h0123]=16'h0256;
      mem0[16'h0124]=16'h0300;
      mem1[16'h0124]=16'hd333;
      mem0[16'h0125]=16'h0170;
      mem1[16'h0125]=16'h000a;
      mem0[16'h0126]=16'h0380;
      mem1[16'h0126]=16'he555;
      mem0[16'h0127]=16'h0160;
      mem1[16'h0127]=16'h0f18;
      mem0[16'h0128]=16'h3650;
      mem1[16'h0128]=16'h0c45;
      mem0[16'h0129]=16'h0160;
      mem1[16'h0129]=16'h0890;
      mem0[16'h012a]=16'h01c0;
      mem1[16'h012a]=16'h0104;
      mem0[16'h012b]=16'h0164;
      mem1[16'h012b]=16'h0a78;
      mem0[16'h012c]=16'h0160;
      mem1[16'h012c]=16'h087c;
      mem0[16'h012d]=16'h01c0;
      mem1[16'h012d]=16'h0114;
      mem0[16'h012e]=16'h3a24;
      mem1[16'h012e]=16'h0104;
      mem0[16'h012f]=16'h0160;
      mem1[16'h012f]=16'h089c;
      mem0[16'h0130]=16'h01c0;
      mem1[16'h0130]=16'h1220;
      mem0[16'h0131]=16'h0160;
      mem1[16'h0131]=16'h0ad4;
      mem0[16'h0132]=16'h01c0;
      mem1[16'h0132]=16'h0160;
      mem0[16'h0133]=16'h0920;
      mem1[16'h0133]=16'h01c0;
      mem0[16'h0134]=16'h0164;
      mem1[16'h0134]=16'h0f00;
      mem0[16'h0135]=16'h0160;
      mem1[16'h0135]=16'h09c2;
      mem0[16'h0136]=16'h01c0;
      mem1[16'h0136]=16'hd222;
      mem0[16'h0137]=16'h0170;
      mem1[16'h0137]=16'h0012;
      mem0[16'h0138]=16'h0380;
      mem1[16'h0138]=16'h0114;
      mem0[16'h0139]=16'h0841;
      mem1[16'h0139]=16'h0160;
      mem0[16'h013a]=16'h0f18;
      mem1[16'h013a]=16'h3440;
      mem0[16'h013b]=16'h0170;
      mem1[16'h013b]=16'hffb4;
      mem0[16'h013c]=16'h01f0;
      mem1[16'h013c]=16'h102d;
      mem0[16'h013d]=16'hf220;
      mem1[16'h013d]=16'h0170;
      mem0[16'h013e]=16'h0012;
      mem1[16'h013e]=16'h0380;
      mem0[16'h013f]=16'h0114;
      mem1[16'h013f]=16'h0941;
      mem0[16'h0140]=16'h0160;
      mem1[16'h0140]=16'h0f18;
      mem0[16'h0141]=16'h3440;
      mem1[16'h0141]=16'h0170;
      mem0[16'h0142]=16'hff9a;
      mem1[16'h0142]=16'h01f0;
      mem0[16'h0143]=16'h102e;
      mem1[16'h0143]=16'hf220;
      mem0[16'h0144]=16'h0170;
      mem1[16'h0144]=16'h0010;
      mem0[16'h0145]=16'h0380;
      mem1[16'h0145]=16'h0114;
      mem0[16'h0146]=16'h0160;
      mem1[16'h0146]=16'h0f18;
      mem0[16'h0147]=16'h3440;
      mem1[16'h0147]=16'h0160;
      mem0[16'h0148]=16'h01fc;
      mem1[16'h0148]=16'h01e0;
      mem0[16'h0149]=16'h0160;
      mem1[16'h0149]=16'h09e6;
      mem0[16'h014a]=16'h01c0;
      mem1[16'h014a]=16'hd333;
      mem0[16'h014b]=16'h0114;
      mem1[16'h014b]=16'h0160;
      mem0[16'h014c]=16'h0256;
      mem1[16'h014c]=16'h0340;
      mem0[16'h014d]=16'h3854;
      mem1[16'h014d]=16'h0841;
      mem0[16'h014e]=16'h0160;
      mem1[16'h014e]=16'h0f18;
      mem0[16'h014f]=16'h3440;
      mem1[16'h014f]=16'h0170;
      mem0[16'h0150]=16'hff62;
      mem1[16'h0150]=16'h01f0;
      mem0[16'h0151]=16'h0841;
      mem1[16'h0151]=16'h0160;
      mem0[16'h0152]=16'h09c2;
      mem1[16'h0152]=16'h01c0;
      mem0[16'h0153]=16'h0160;
      mem1[16'h0153]=16'h09e6;
      mem0[16'h0154]=16'h01c0;
      mem1[16'h0154]=16'h0160;
      mem0[16'h0155]=16'h09c2;
      mem1[16'h0155]=16'h01c0;
      mem0[16'h0156]=16'hd222;
      mem1[16'h0156]=16'h0160;
      mem0[16'h0157]=16'h0256;
      mem1[16'h0157]=16'h0300;
      mem0[16'h0158]=16'hd333;
      mem1[16'h0158]=16'h0170;
      mem0[16'h0159]=16'h0004;
      mem1[16'h0159]=16'h0380;
      mem0[16'h015a]=16'h1500;
      mem1[16'h015a]=16'h0160;
      mem0[16'h015b]=16'h0ab8;
      mem1[16'h015b]=16'h01c0;
      mem0[16'h015c]=16'h0160;
      mem1[16'h015c]=16'h09d4;
      mem0[16'h015d]=16'h01c0;
      mem1[16'h015d]=16'h1053;
      mem0[16'h015e]=16'hf220;
      mem1[16'h015e]=16'h0170;
      mem0[16'h015f]=16'h00c0;
      mem1[16'h015f]=16'h03c0;
      mem0[16'h0160]=16'h103a;
      mem1[16'h0160]=16'hf220;
      mem0[16'h0161]=16'h0170;
      mem1[16'h0161]=16'h0022;
      mem0[16'h0162]=16'h03c0;
      mem1[16'h0162]=16'h100d;
      mem0[16'h0163]=16'hf220;
      mem1[16'h0163]=16'h0170;
      mem0[16'h0164]=16'hffd8;
      mem1[16'h0164]=16'h03c0;
      mem0[16'h0165]=16'h100a;
      mem1[16'h0165]=16'hf220;
      mem0[16'h0166]=16'h0170;
      mem1[16'h0166]=16'hffce;
      mem0[16'h0167]=16'h03c0;
      mem1[16'h0167]=16'h0160;
      mem0[16'h0168]=16'h0ab8;
      mem1[16'h0168]=16'h01c0;
      mem0[16'h0169]=16'h0170;
      mem1[16'h0169]=16'hffe2;
      mem0[16'h016a]=16'h01f0;
      mem1[16'h016a]=16'h0160;
      mem0[16'h016b]=16'h08c2;
      mem1[16'h016b]=16'h01c0;
      mem0[16'h016c]=16'h3c29;
      mem1[16'h016c]=16'h3c28;
      mem0[16'h016d]=16'h0160;
      mem1[16'h016d]=16'h08c2;
      mem0[16'h016e]=16'h01c0;
      mem1[16'h016e]=16'h8992;
      mem0[16'h016f]=16'h0628;
      mem1[16'h016f]=16'h3c24;
      mem0[16'h0170]=16'h0160;
      mem1[16'h0170]=16'h08c2;
      mem0[16'h0171]=16'h01c0;
      mem1[16'h0171]=16'hd442;
      mem0[16'h0172]=16'h8992;
      mem1[16'h0172]=16'h8445;
      mem0[16'h0173]=16'h0160;
      mem1[16'h0173]=16'h08c2;
      mem0[16'h0174]=16'h01c0;
      mem1[16'h0174]=16'h0160;
      mem0[16'h0175]=16'h0f1b;
      mem1[16'h0175]=16'h3820;
      mem0[16'h0176]=16'h8992;
      mem1[16'h0176]=16'hd888;
      mem0[16'h0177]=16'h0170;
      mem1[16'h0177]=16'h0024;
      mem0[16'h0178]=16'h03c0;
      mem1[16'h0178]=16'h0160;
      mem0[16'h0179]=16'h08c2;
      mem1[16'h0179]=16'h01c0;
      mem0[16'h017a]=16'h8992;
      mem1[16'h017a]=16'he666;
      mem0[16'h017b]=16'h0160;
      mem1[16'h017b]=16'h0f1b;
      mem0[16'h017c]=16'h3a60;
      mem1[16'h017c]=16'hd666;
      mem0[16'h017d]=16'h0170;
      mem1[16'h017d]=16'h0006;
      mem0[16'h017e]=16'h0380;
      mem1[16'h017e]=16'h3824;
      mem0[16'h017f]=16'h0841;
      mem1[16'h017f]=16'h0170;
      mem0[16'h0180]=16'hffe0;
      mem1[16'h0180]=16'h0a80;
      mem0[16'h0181]=16'h0160;
      mem1[16'h0181]=16'h08c2;
      mem0[16'h0182]=16'h01c0;
      mem1[16'h0182]=16'h8992;
      mem0[16'h0183]=16'h10ff;
      mem1[16'h0183]=16'hc990;
      mem0[16'h0184]=16'hd999;
      mem1[16'h0184]=16'h0170;
      mem0[16'h0185]=16'h0018;
      mem1[16'h0185]=16'h0380;
      mem0[16'h0186]=16'he666;
      mem1[16'h0186]=16'h0160;
      mem0[16'h0187]=16'h0f1b;
      mem1[16'h0187]=16'h3a60;
      mem0[16'h0188]=16'hd666;
      mem1[16'h0188]=16'h0160;
      mem0[16'h0189]=16'h059e;
      mem1[16'h0189]=16'h0340;
      mem0[16'h018a]=16'h0160;
      mem1[16'h018a]=16'h01fc;
      mem0[16'h018b]=16'h01e0;
      mem1[16'h018b]=16'h0164;
      mem0[16'h018c]=16'h0a53;
      mem1[16'h018c]=16'h0160;
      mem0[16'h018d]=16'h087c;
      mem1[16'h018d]=16'h01c0;
      mem0[16'h018e]=16'h0160;
      mem1[16'h018e]=16'h01fc;
      mem0[16'h018f]=16'h01e0;
      mem1[16'h018f]=16'h0160;
      mem0[16'h0190]=16'h0ab8;
      mem1[16'h0190]=16'h01c0;
      mem0[16'h0191]=16'h0160;
      mem1[16'h0191]=16'h0f1b;
      mem0[16'h0192]=16'h3820;
      mem1[16'h0192]=16'h0160;
      mem0[16'h0193]=16'h08c2;
      mem1[16'h0193]=16'h01c0;
      mem0[16'h0194]=16'h3c28;
      mem1[16'h0194]=16'h3c29;
      mem0[16'h0195]=16'h0160;
      mem1[16'h0195]=16'h08c2;
      mem0[16'h0196]=16'h01c0;
      mem1[16'h0196]=16'h8992;
      mem0[16'h0197]=16'h0628;
      mem1[16'h0197]=16'h3c24;
      mem0[16'h0198]=16'h0160;
      mem1[16'h0198]=16'h08c2;
      mem0[16'h0199]=16'h01c0;
      mem1[16'h0199]=16'hd442;
      mem0[16'h019a]=16'h8992;
      mem1[16'h019a]=16'h8445;
      mem0[16'h019b]=16'h0983;
      mem1[16'h019b]=16'h0170;
      mem0[16'h019c]=16'h0026;
      mem1[16'h019c]=16'h03c0;
      mem0[16'h019d]=16'h0160;
      mem1[16'h019d]=16'h08c2;
      mem0[16'h019e]=16'h01c0;
      mem1[16'h019e]=16'h8992;
      mem0[16'h019f]=16'he666;
      mem1[16'h019f]=16'h0160;
      mem0[16'h01a0]=16'h0f1b;
      mem1[16'h01a0]=16'h3a60;
      mem0[16'h01a1]=16'h1031;
      mem1[16'h01a1]=16'hf660;
      mem0[16'h01a2]=16'h0170;
      mem1[16'h01a2]=16'h0006;
      mem0[16'h01a3]=16'h0380;
      mem1[16'h01a3]=16'h3824;
      mem0[16'h01a4]=16'h0841;
      mem1[16'h01a4]=16'h0170;
      mem0[16'h01a5]=16'hffde;
      mem1[16'h01a5]=16'h0a80;
      mem0[16'h01a6]=16'h0160;
      mem1[16'h01a6]=16'h08c2;
      mem0[16'h01a7]=16'h01c0;
      mem1[16'h01a7]=16'h8992;
      mem0[16'h01a8]=16'h10ff;
      mem1[16'h01a8]=16'hc990;
      mem0[16'h01a9]=16'h10ff;
      mem1[16'h01a9]=16'hf990;
      mem0[16'h01aa]=16'h0170;
      mem1[16'h01aa]=16'h002e;
      mem0[16'h01ab]=16'h0380;
      mem1[16'h01ab]=16'he666;
      mem0[16'h01ac]=16'h0160;
      mem1[16'h01ac]=16'h0f1b;
      mem0[16'h01ad]=16'h3a60;
      mem1[16'h01ad]=16'h1037;
      mem0[16'h01ae]=16'hf660;
      mem1[16'h01ae]=16'h0170;
      mem0[16'h01af]=16'h0026;
      mem1[16'h01af]=16'h03c0;
      mem0[16'h01b0]=16'h1038;
      mem1[16'h01b0]=16'hf660;
      mem0[16'h01b1]=16'h0170;
      mem1[16'h01b1]=16'h001c;
      mem0[16'h01b2]=16'h03c0;
      mem1[16'h01b2]=16'h1039;
      mem0[16'h01b3]=16'hf660;
      mem1[16'h01b3]=16'h0170;
      mem0[16'h01b4]=16'h0012;
      mem1[16'h01b4]=16'h03c0;
      mem0[16'h01b5]=16'h0160;
      mem1[16'h01b5]=16'h059e;
      mem0[16'h01b6]=16'h01e0;
      mem1[16'h01b6]=16'h0164;
      mem0[16'h01b7]=16'h0a60;
      mem1[16'h01b7]=16'h0160;
      mem0[16'h01b8]=16'h087c;
      mem1[16'h01b8]=16'h01c0;
      mem0[16'h01b9]=16'h0160;
      mem1[16'h01b9]=16'h01fc;
      mem0[16'h01ba]=16'h01e0;
      mem1[16'h01ba]=16'h0841;
      mem0[16'h01bb]=16'he222;
      mem1[16'h01bb]=16'h3a24;
      mem0[16'h01bc]=16'h0160;
      mem1[16'h01bc]=16'h09d4;
      mem0[16'h01bd]=16'h01c0;
      mem1[16'h01bd]=16'h1049;
      mem0[16'h01be]=16'hf220;
      mem1[16'h01be]=16'h0170;
      mem0[16'h01bf]=16'h000c;
      mem1[16'h01bf]=16'h03c0;
      mem0[16'h01c0]=16'h1053;
      mem1[16'h01c0]=16'hf220;
      mem0[16'h01c1]=16'h0170;
      mem1[16'h01c1]=16'h000a;
      mem0[16'h01c2]=16'h0380;
      mem1[16'h01c2]=16'h0841;
      mem0[16'h01c3]=16'h0160;
      mem1[16'h01c3]=16'h0f1a;
      mem0[16'h01c4]=16'h3820;
      mem1[16'h01c4]=16'h0160;
      mem0[16'h01c5]=16'h09c2;
      mem1[16'h01c5]=16'h01c0;
      mem0[16'h01c6]=16'h0160;
      mem1[16'h01c6]=16'h09e6;
      mem0[16'h01c7]=16'h01c0;
      mem1[16'h01c7]=16'hd333;
      mem0[16'h01c8]=16'h0170;
      mem1[16'h01c8]=16'h0038;
      mem0[16'h01c9]=16'h03c0;
      mem1[16'h01c9]=16'h3c58;
      mem0[16'h01ca]=16'h0160;
      mem1[16'h01ca]=16'h09c2;
      mem0[16'h01cb]=16'h01c0;
      mem1[16'h01cb]=16'h102c;
      mem0[16'h01cc]=16'hf220;
      mem1[16'h01cc]=16'h0170;
      mem0[16'h01cd]=16'h0026;
      mem1[16'h01cd]=16'h0380;
      mem0[16'h01ce]=16'h0841;
      mem1[16'h01ce]=16'h0160;
      mem0[16'h01cf]=16'h09c2;
      mem1[16'h01cf]=16'h01c0;
      mem0[16'h01d0]=16'h0160;
      mem1[16'h01d0]=16'h09e6;
      mem0[16'h01d1]=16'h01c0;
      mem1[16'h01d1]=16'hd333;
      mem0[16'h01d2]=16'h0170;
      mem1[16'h01d2]=16'h0010;
      mem0[16'h01d3]=16'h03c0;
      mem1[16'h01d3]=16'h0160;
      mem0[16'h01d4]=16'h09c2;
      mem1[16'h01d4]=16'h01c0;
      mem0[16'h01d5]=16'hd222;
      mem1[16'h01d5]=16'h0170;
      mem0[16'h01d6]=16'h0008;
      mem1[16'h01d6]=16'h03c0;
      mem0[16'h01d7]=16'h0160;
      mem1[16'h01d7]=16'h0256;
      mem0[16'h01d8]=16'h01e0;
      mem1[16'h01d8]=16'h3c84;
      mem0[16'h01d9]=16'h0c45;
      mem1[16'h01d9]=16'h0841;
      mem0[16'h01da]=16'h9445;
      mem1[16'h01da]=16'h0160;
      mem0[16'h01db]=16'h07aa;
      mem1[16'h01db]=16'h01c0;
      mem0[16'h01dc]=16'hd444;
      mem1[16'h01dc]=16'h0170;
      mem0[16'h01dd]=16'hfff4;
      mem1[16'h01dd]=16'h0380;
      mem0[16'h01de]=16'he666;
      mem1[16'h01de]=16'h0160;
      mem0[16'h01df]=16'h0f1a;
      mem1[16'h01df]=16'h3a60;
      mem0[16'h01e0]=16'h1049;
      mem1[16'h01e0]=16'hf660;
      mem0[16'h01e1]=16'h0170;
      mem1[16'h01e1]=16'h0012;
      mem0[16'h01e2]=16'h0380;
      mem1[16'h01e2]=16'h0164;
      mem0[16'h01e3]=16'h0a7c;
      mem1[16'h01e3]=16'h0160;
      mem0[16'h01e4]=16'h087c;
      mem1[16'h01e4]=16'h01c0;
      mem0[16'h01e5]=16'h0160;
      mem1[16'h01e5]=16'h01fc;
      mem0[16'h01e6]=16'h01e0;
      mem1[16'h01e6]=16'h0164;
      mem0[16'h01e7]=16'h0a8a;
      mem1[16'h01e7]=16'h0160;
      mem0[16'h01e8]=16'h087c;
      mem1[16'h01e8]=16'h01c0;
      mem0[16'h01e9]=16'h0160;
      mem1[16'h01e9]=16'h01fc;
      mem0[16'h01ea]=16'h01e0;
      mem1[16'h01ea]=16'h1810;
      mem0[16'h01eb]=16'hf448;
      mem1[16'h01eb]=16'h0170;
      mem0[16'h01ec]=16'h0004;
      mem1[16'h01ec]=16'h0390;
      mem0[16'h01ed]=16'h3c48;
      mem1[16'h01ed]=16'h9448;
      mem0[16'h01ee]=16'he666;
      mem1[16'h01ee]=16'h0160;
      mem0[16'h01ef]=16'h0f1a;
      mem1[16'h01ef]=16'h3a60;
      mem0[16'h01f0]=16'h1049;
      mem1[16'h01f0]=16'hf660;
      mem0[16'h01f1]=16'h0170;
      mem1[16'h01f1]=16'h005a;
      mem0[16'h01f2]=16'h0380;
      mem1[16'h01f2]=16'h123a;
      mem0[16'h01f3]=16'h0160;
      mem1[16'h01f3]=16'h0ad4;
      mem0[16'h01f4]=16'h01c0;
      mem1[16'h01f4]=16'h3c82;
      mem0[16'h01f5]=16'h0160;
      mem1[16'h01f5]=16'h089c;
      mem0[16'h01f6]=16'h01c0;
      mem1[16'h01f6]=16'h3c89;
      mem0[16'h01f7]=16'h3c52;
      mem1[16'h01f7]=16'h0528;
      mem0[16'h01f8]=16'h8992;
      mem1[16'h01f8]=16'h0160;
      mem0[16'h01f9]=16'h089c;
      mem1[16'h01f9]=16'h01c0;
      mem0[16'h01fa]=16'hc225;
      mem1[16'h01fa]=16'h10ff;
      mem0[16'h01fb]=16'hc220;
      mem1[16'h01fb]=16'h8992;
      mem0[16'h01fc]=16'h0160;
      mem1[16'h01fc]=16'h089c;
      mem0[16'h01fd]=16'h01c0;
      mem1[16'h01fd]=16'he222;
      mem0[16'h01fe]=16'h0160;
      mem1[16'h01fe]=16'h089c;
      mem0[16'h01ff]=16'h01c0;
      mem1[16'h01ff]=16'he222;
      mem0[16'h0200]=16'h3a25;
      mem1[16'h0200]=16'h8992;
      mem0[16'h0201]=16'h0160;
      mem1[16'h0201]=16'h089c;
      mem0[16'h0202]=16'h01c0;
      mem1[16'h0202]=16'h0851;
      mem0[16'h0203]=16'h0170;
      mem1[16'h0203]=16'hffee;
      mem0[16'h0204]=16'h0a80;
      mem1[16'h0204]=16'h0159;
      mem0[16'h0205]=16'h3c92;
      mem1[16'h0205]=16'h0160;
      mem0[16'h0206]=16'h089c;
      mem1[16'h0206]=16'h01c0;
      mem0[16'h0207]=16'h0160;
      mem1[16'h0207]=16'h0910;
      mem0[16'h0208]=16'h01e0;
      mem1[16'h0208]=16'h1253;
      mem0[16'h0209]=16'h0160;
      mem1[16'h0209]=16'h0ad4;
      mem0[16'h020a]=16'h01c0;
      mem1[16'h020a]=16'h1231;
      mem0[16'h020b]=16'h0160;
      mem1[16'h020b]=16'h0ad4;
      mem0[16'h020c]=16'h01c0;
      mem1[16'h020c]=16'h0883;
      mem0[16'h020d]=16'h3c89;
      mem1[16'h020d]=16'h3c82;
      mem0[16'h020e]=16'h0160;
      mem1[16'h020e]=16'h089c;
      mem0[16'h020f]=16'h01c0;
      mem1[16'h020f]=16'h3c42;
      mem0[16'h0210]=16'h0528;
      mem1[16'h0210]=16'h3c29;
      mem0[16'h0211]=16'h0160;
      mem1[16'h0211]=16'h089c;
      mem0[16'h0212]=16'h01c0;
      mem1[16'h0212]=16'h3c42;
      mem0[16'h0213]=16'h10ff;
      mem1[16'h0213]=16'hc220;
      mem0[16'h0214]=16'h3c29;
      mem1[16'h0214]=16'h0160;
      mem0[16'h0215]=16'h089c;
      mem1[16'h0215]=16'h01c0;
      mem0[16'h0216]=16'he222;
      mem1[16'h0216]=16'h3a25;
      mem0[16'h0217]=16'h8992;
      mem1[16'h0217]=16'h0160;
      mem0[16'h0218]=16'h089c;
      mem1[16'h0218]=16'h01c0;
      mem0[16'h0219]=16'h0851;
      mem1[16'h0219]=16'h0170;
      mem0[16'h021a]=16'hffee;
      mem1[16'h021a]=16'h0a80;
      mem0[16'h021b]=16'h0149;
      mem1[16'h021b]=16'h3c92;
      mem0[16'h021c]=16'h0160;
      mem1[16'h021c]=16'h089c;
      mem0[16'h021d]=16'h01c0;
      mem1[16'h021d]=16'h0160;
      mem0[16'h021e]=16'h0910;
      mem1[16'h021e]=16'h01e0;
      mem0[16'h021f]=16'h3a24;
      mem1[16'h021f]=16'hc222;
      mem0[16'h0220]=16'h0084;
      mem1[16'h0220]=16'h0160;
      mem0[16'h0221]=16'h0ad4;
      mem1[16'h0221]=16'h01c0;
      mem0[16'h0222]=16'h0841;
      mem1[16'h0222]=16'h0170;
      mem0[16'h0223]=16'hffee;
      mem1[16'h0223]=16'h01f0;
      mem0[16'h0224]=16'h3c42;
      mem1[16'h0224]=16'h0428;
      mem0[16'h0225]=16'h0160;
      mem1[16'h0225]=16'h089c;
      mem0[16'h0226]=16'h01c0;
      mem1[16'h0226]=16'h3c42;
      mem0[16'h0227]=16'h3c26;
      mem1[16'h0227]=16'h0424;
      mem0[16'h0228]=16'h0160;
      mem1[16'h0228]=16'h08a8;
      mem0[16'h0229]=16'h01c0;
      mem1[16'h0229]=16'h3c62;
      mem0[16'h022a]=16'h100f;
      mem1[16'h022a]=16'hc220;
      mem0[16'h022b]=16'h1030;
      mem1[16'h022b]=16'h8220;
      mem0[16'h022c]=16'h103a;
      mem1[16'h022c]=16'hf220;
      mem0[16'h022d]=16'h0160;
      mem1[16'h022d]=16'h0ad4;
      mem0[16'h022e]=16'h0350;
      mem1[16'h022e]=16'h0827;
      mem0[16'h022f]=16'h0160;
      mem1[16'h022f]=16'h0ad4;
      mem0[16'h0230]=16'h01e0;
      mem1[16'h0230]=16'he222;
      mem0[16'h0231]=16'h0160;
      mem1[16'h0231]=16'h08cc;
      mem0[16'h0232]=16'h01c0;
      mem1[16'h0232]=16'h0624;
      mem0[16'h0233]=16'h0108;
      mem1[16'h0233]=16'h3c28;
      mem0[16'h0234]=16'h0160;
      mem1[16'h0234]=16'h0ab8;
      mem0[16'h0235]=16'h01c0;
      mem1[16'h0235]=16'h0160;
      mem0[16'h0236]=16'h09d4;
      mem1[16'h0236]=16'h01c0;
      mem0[16'h0237]=16'h1030;
      mem1[16'h0237]=16'hf220;
      mem0[16'h0238]=16'h0170;
      mem1[16'h0238]=16'h0028;
      mem0[16'h0239]=16'h03d0;
      mem1[16'h0239]=16'h103a;
      mem0[16'h023a]=16'hf220;
      mem1[16'h023a]=16'h0170;
      mem0[16'h023b]=16'h0018;
      mem1[16'h023b]=16'h03d0;
      mem0[16'h023c]=16'h1041;
      mem1[16'h023c]=16'hf220;
      mem0[16'h023d]=16'h0170;
      mem1[16'h023d]=16'h0014;
      mem0[16'h023e]=16'h03d0;
      mem1[16'h023e]=16'h1047;
      mem0[16'h023f]=16'hf220;
      mem1[16'h023f]=16'h0170;
      mem0[16'h0240]=16'h000a;
      mem1[16'h0240]=16'h0390;
      mem0[16'h0241]=16'h0927;
      mem1[16'h0241]=16'h1030;
      mem0[16'h0242]=16'h9220;
      mem1[16'h0242]=16'hd228;
      mem0[16'h0243]=16'h0118;
      mem1[16'h0243]=16'h0002;
      mem0[16'h0244]=16'h120d;
      mem1[16'h0244]=16'h0160;
      mem0[16'h0245]=16'h0ad4;
      mem1[16'h0245]=16'h01c0;
      mem0[16'h0246]=16'h120a;
      mem1[16'h0246]=16'h0160;
      mem0[16'h0247]=16'h0ad4;
      mem1[16'h0247]=16'h01e0;
      mem0[16'h0248]=16'h010a;
      mem1[16'h0248]=16'h0108;
      mem0[16'h0249]=16'h016a;
      mem1[16'h0249]=16'h0f00;
      mem0[16'h024a]=16'h1800;
      mem1[16'h024a]=16'h0160;
      mem0[16'h024b]=16'h0ab8;
      mem1[16'h024b]=16'h01c0;
      mem0[16'h024c]=16'h100d;
      mem1[16'h024c]=16'hf220;
      mem0[16'h024d]=16'h0170;
      mem1[16'h024d]=16'h007a;
      mem0[16'h024e]=16'h03c0;
      mem1[16'h024e]=16'h100a;
      mem0[16'h024f]=16'hf220;
      mem1[16'h024f]=16'h0170;
      mem0[16'h0250]=16'h0070;
      mem1[16'h0250]=16'h03c0;
      mem0[16'h0251]=16'h1008;
      mem1[16'h0251]=16'hf220;
      mem0[16'h0252]=16'h0170;
      mem1[16'h0252]=16'h003c;
      mem0[16'h0253]=16'h03c0;
      mem1[16'h0253]=16'h107f;
      mem0[16'h0254]=16'hf220;
      mem1[16'h0254]=16'h0170;
      mem0[16'h0255]=16'h0032;
      mem1[16'h0255]=16'h03c0;
      mem0[16'h0256]=16'h1020;
      mem1[16'h0256]=16'hf220;
      mem0[16'h0257]=16'h0170;
      mem1[16'h0257]=16'hffca;
      mem0[16'h0258]=16'h03d0;
      mem1[16'h0258]=16'h1080;
      mem0[16'h0259]=16'hf220;
      mem1[16'h0259]=16'h0170;
      mem0[16'h025a]=16'hffc0;
      mem1[16'h025a]=16'h0390;
      mem0[16'h025b]=16'h100f;
      mem1[16'h025b]=16'hf880;
      mem0[16'h025c]=16'h0170;
      mem1[16'h025c]=16'hffb6;
      mem0[16'h025d]=16'h0390;
      mem1[16'h025d]=16'h0881;
      mem0[16'h025e]=16'h0160;
      mem1[16'h025e]=16'h0ad4;
      mem0[16'h025f]=16'h01c0;
      mem1[16'h025f]=16'h382a;
      mem0[16'h0260]=16'h08a1;
      mem1[16'h0260]=16'h0170;
      mem0[16'h0261]=16'hffa4;
      mem1[16'h0261]=16'h01f0;
      mem0[16'h0262]=16'hc888;
      mem1[16'h0262]=16'h0170;
      mem0[16'h0263]=16'hff9c;
      mem1[16'h0263]=16'h03c0;
      mem0[16'h0264]=16'h0981;
      mem1[16'h0264]=16'h09a1;
      mem0[16'h0265]=16'h1208;
      mem1[16'h0265]=16'h0160;
      mem0[16'h0266]=16'h0ad4;
      mem1[16'h0266]=16'h01c0;
      mem0[16'h0267]=16'h1220;
      mem1[16'h0267]=16'h0160;
      mem0[16'h0268]=16'h0ad4;
      mem1[16'h0268]=16'h01c0;
      mem0[16'h0269]=16'h1208;
      mem1[16'h0269]=16'h0160;
      mem0[16'h026a]=16'h0ad4;
      mem1[16'h026a]=16'h01c0;
      mem0[16'h026b]=16'h0170;
      mem1[16'h026b]=16'hff7a;
      mem0[16'h026c]=16'h01f0;
      mem1[16'h026c]=16'h0160;
      mem0[16'h026d]=16'h0910;
      mem1[16'h026d]=16'h01c0;
      mem0[16'h026e]=16'h1000;
      mem1[16'h026e]=16'h380a;
      mem0[16'h026f]=16'h0118;
      mem1[16'h026f]=16'h011a;
      mem0[16'h0270]=16'h0002;
      mem1[16'h0270]=16'he222;
      mem0[16'h0271]=16'h3a24;
      mem1[16'h0271]=16'h1020;
      mem0[16'h0272]=16'hf220;
      mem1[16'h0272]=16'h0080;
      mem0[16'h0273]=16'h0841;
      mem1[16'h0273]=16'h0170;
      mem0[16'h0274]=16'hfff0;
      mem1[16'h0274]=16'h01f0;
      mem0[16'h0275]=16'h1061;
      mem1[16'h0275]=16'hf220;
      mem0[16'h0276]=16'h0085;
      mem1[16'h0276]=16'h107b;
      mem0[16'h0277]=16'hf220;
      mem1[16'h0277]=16'h0081;
      mem0[16'h0278]=16'h20e0;
      mem1[16'h0278]=16'h8220;
      mem0[16'h0279]=16'h0002;
      mem1[16'h0279]=16'he555;
      mem0[16'h027a]=16'he333;
      mem1[16'h027a]=16'he222;
      mem0[16'h027b]=16'h3a24;
      mem1[16'h027b]=16'h0160;
      mem0[16'h027c]=16'h09d4;
      mem1[16'h027c]=16'h01c0;
      mem0[16'h027d]=16'h1030;
      mem1[16'h027d]=16'hf220;
      mem0[16'h027e]=16'h0170;
      mem1[16'h027e]=16'h0034;
      mem0[16'h027f]=16'h03d0;
      mem1[16'h027f]=16'h103a;
      mem0[16'h0280]=16'hf220;
      mem1[16'h0280]=16'h0170;
      mem0[16'h0281]=16'h0018;
      mem1[16'h0281]=16'h03d0;
      mem0[16'h0282]=16'h1041;
      mem1[16'h0282]=16'hf220;
      mem0[16'h0283]=16'h0170;
      mem1[16'h0283]=16'h0020;
      mem0[16'h0284]=16'h03d0;
      mem1[16'h0284]=16'h1047;
      mem0[16'h0285]=16'hf220;
      mem1[16'h0285]=16'h0170;
      mem0[16'h0286]=16'h0016;
      mem1[16'h0286]=16'h0390;
      mem0[16'h0287]=16'h0927;
      mem1[16'h0287]=16'h1030;
      mem0[16'h0288]=16'h9220;
      mem1[16'h0288]=16'h0654;
      mem0[16'h0289]=16'hd552;
      mem1[16'h0289]=16'h0841;
      mem0[16'h028a]=16'h0831;
      mem1[16'h028a]=16'h0170;
      mem0[16'h028b]=16'hffbc;
      mem1[16'h028b]=16'h01f0;
      mem0[16'h028c]=16'h0002;
      mem1[16'h028c]=16'h0002;
      mem0[16'h028d]=16'h0002;
      mem1[16'h028d]=16'h0a0d;
      mem0[16'h028e]=16'h6e55;
      mem1[16'h028e]=16'h7669;
      mem0[16'h028f]=16'h7265;
      mem1[16'h028f]=16'h6173;
      mem0[16'h0290]=16'h206c;
      mem1[16'h0290]=16'h6f4d;
      mem0[16'h0291]=16'h696e;
      mem1[16'h0291]=16'h6f74;
      mem0[16'h0292]=16'h2072;
      mem1[16'h0292]=16'h3848;
      mem0[16'h0293]=16'h0d30;
      mem1[16'h0293]=16'h000a;
      mem0[16'h0294]=16'h205d;
      mem1[16'h0294]=16'h4500;
      mem0[16'h0295]=16'h7272;
      mem1[16'h0295]=16'h726f;
      mem0[16'h0296]=16'h6920;
      mem1[16'h0296]=16'h6568;
      mem0[16'h0297]=16'h0d78;
      mem1[16'h0297]=16'h000a;
      mem0[16'h0298]=16'h7245;
      mem1[16'h0298]=16'h6f72;
      mem0[16'h0299]=16'h2072;
      mem1[16'h0299]=16'h7273;
      mem0[16'h029a]=16'h6365;
      mem1[16'h029a]=16'h0a0d;
      mem0[16'h029b]=16'h4500;
      mem1[16'h029b]=16'h7272;
      mem0[16'h029c]=16'h726f;
      mem1[16'h029c]=16'h0a0d;
      mem0[16'h029d]=16'h2000;
      mem1[16'h029d]=16'h003a;
      mem0[16'h029e]=16'h3a20;
      mem1[16'h029e]=16'h0020;
      mem0[16'h029f]=16'h303a;
      mem1[16'h029f]=16'h3030;
      mem0[16'h02a0]=16'h3030;
      mem1[16'h02a0]=16'h3030;
      mem0[16'h02a1]=16'h4631;
      mem1[16'h02a1]=16'h0d46;
      mem0[16'h02a2]=16'h000a;
      mem1[16'h02a2]=16'h3953;
      mem0[16'h02a3]=16'h3330;
      mem1[16'h02a3]=16'h3030;
      mem0[16'h02a4]=16'h3030;
      mem1[16'h02a4]=16'h4346;
      mem0[16'h02a5]=16'h0a0d;
      mem1[16'h02a5]=16'h4800;
      mem0[16'h02a6]=16'h3038;
      mem1[16'h02a6]=16'h3128;
      mem0[16'h02a7]=16'h2936;
      mem1[16'h02a7]=16'h0a0d;
      mem0[16'h02a8]=16'h4800;
      mem1[16'h02a8]=16'h3038;
      mem0[16'h02a9]=16'h3328;
      mem1[16'h02a9]=16'h2932;
      mem0[16'h02aa]=16'h0a0d;
      mem1[16'h02aa]=16'h5200;
      mem0[16'h02ab]=16'h5453;
      mem1[16'h02ab]=16'h3320;
      mem0[16'h02ac]=16'h4838;
      mem1[16'h02ac]=16'h0a0d;
      mem0[16'h02ad]=16'hff00;
      mem1[16'h02ad]=16'h0002;
      mem0[16'h02ae]=16'h0160;
      mem1[16'h02ae]=16'h0aca;
      mem0[16'h02af]=16'h01c0;
      mem1[16'h02af]=16'h0170;
      mem0[16'h02b0]=16'hfff6;
      mem1[16'h02b0]=16'h03c0;
      mem0[16'h02b1]=16'h1000;
      mem1[16'h02b1]=16'h3b20;
      mem0[16'h02b2]=16'h0002;
      mem1[16'h02b2]=16'he222;
      mem0[16'h02b3]=16'h1001;
      mem1[16'h02b3]=16'h3b20;
      mem0[16'h02b4]=16'hd222;
      mem1[16'h02b4]=16'h0002;
      mem0[16'h02b5]=16'h1000;
      mem1[16'h02b5]=16'h3920;
      mem0[16'h02b6]=16'h0002;
      mem1[16'h02b6]=16'hffff;
      mem0[16'h02b7]=16'hffff;
      mem1[16'h02b7]=16'hffff;
      mem0[16'h02b8]=16'hffff;
      mem1[16'h02b8]=16'hffff;
      mem0[16'h02b9]=16'hffff;
      mem1[16'h02b9]=16'hffff;
      mem0[16'h02ba]=16'hffff;
      mem1[16'h02ba]=16'hffff;
      mem0[16'h02bb]=16'hffff;
      mem1[16'h02bb]=16'hffff;
      mem0[16'h02bc]=16'hffff;
      mem1[16'h02bc]=16'hffff;
      mem0[16'h02bd]=16'hffff;
      mem1[16'h02bd]=16'hffff;
      mem0[16'h02be]=16'hffff;
      mem1[16'h02be]=16'hffff;
      mem0[16'h02bf]=16'hffff;
      mem1[16'h02bf]=16'hffff;
      mem0[16'h02c0]=16'hffff;
      mem1[16'h02c0]=16'hffff;
      mem0[16'h02c1]=16'hffff;
      mem1[16'h02c1]=16'hffff;
      mem0[16'h02c2]=16'hffff;
      mem1[16'h02c2]=16'hffff;
      mem0[16'h02c3]=16'hffff;
      mem1[16'h02c3]=16'hffff;
      mem0[16'h02c4]=16'hffff;
      mem1[16'h02c4]=16'hffff;
      mem0[16'h02c5]=16'hffff;
      mem1[16'h02c5]=16'hffff;
      mem0[16'h02c6]=16'hffff;
      mem1[16'h02c6]=16'hffff;
      mem0[16'h02c7]=16'hffff;
      mem1[16'h02c7]=16'hffff;
      mem0[16'h02c8]=16'hffff;
      mem1[16'h02c8]=16'hffff;
      mem0[16'h02c9]=16'hffff;
      mem1[16'h02c9]=16'hffff;
      mem0[16'h02ca]=16'hffff;
      mem1[16'h02ca]=16'hffff;
      mem0[16'h02cb]=16'hffff;
      mem1[16'h02cb]=16'hffff;
      mem0[16'h02cc]=16'hffff;
      mem1[16'h02cc]=16'hffff;
      mem0[16'h02cd]=16'hffff;
      mem1[16'h02cd]=16'hffff;
      mem0[16'h02ce]=16'hffff;
      mem1[16'h02ce]=16'hffff;
      mem0[16'h02cf]=16'hffff;
      mem1[16'h02cf]=16'hffff;
      mem0[16'h02d0]=16'hffff;
      mem1[16'h02d0]=16'hffff;
      mem0[16'h02d1]=16'hffff;
      mem1[16'h02d1]=16'hffff;
      mem0[16'h02d2]=16'hffff;
      mem1[16'h02d2]=16'hffff;
      mem0[16'h02d3]=16'hffff;
      mem1[16'h02d3]=16'hffff;
      mem0[16'h02d4]=16'hffff;
      mem1[16'h02d4]=16'hffff;
      mem0[16'h02d5]=16'hffff;
      mem1[16'h02d5]=16'hffff;
      mem0[16'h02d6]=16'hffff;
      mem1[16'h02d6]=16'hffff;
      mem0[16'h02d7]=16'hffff;
      mem1[16'h02d7]=16'hffff;
      mem0[16'h02d8]=16'hffff;
      mem1[16'h02d8]=16'hffff;
      mem0[16'h02d9]=16'hffff;
      mem1[16'h02d9]=16'hffff;
      mem0[16'h02da]=16'hffff;
      mem1[16'h02da]=16'hffff;
      mem0[16'h02db]=16'hffff;
      mem1[16'h02db]=16'hffff;
      mem0[16'h02dc]=16'hffff;
      mem1[16'h02dc]=16'hffff;
      mem0[16'h02dd]=16'hffff;
      mem1[16'h02dd]=16'hffff;
      mem0[16'h02de]=16'hffff;
      mem1[16'h02de]=16'hffff;
      mem0[16'h02df]=16'hffff;
      mem1[16'h02df]=16'hffff;
      mem0[16'h02e0]=16'hffff;
      mem1[16'h02e0]=16'hffff;
      mem0[16'h02e1]=16'hffff;
      mem1[16'h02e1]=16'hffff;
      mem0[16'h02e2]=16'hffff;
      mem1[16'h02e2]=16'hffff;
      mem0[16'h02e3]=16'hffff;
      mem1[16'h02e3]=16'hffff;
      mem0[16'h02e4]=16'hffff;
      mem1[16'h02e4]=16'hffff;
      mem0[16'h02e5]=16'hffff;
      mem1[16'h02e5]=16'hffff;
      mem0[16'h02e6]=16'hffff;
      mem1[16'h02e6]=16'hffff;
      mem0[16'h02e7]=16'hffff;
      mem1[16'h02e7]=16'hffff;
      mem0[16'h02e8]=16'hffff;
      mem1[16'h02e8]=16'hffff;
      mem0[16'h02e9]=16'hffff;
      mem1[16'h02e9]=16'hffff;
      mem0[16'h02ea]=16'hffff;
      mem1[16'h02ea]=16'hffff;
      mem0[16'h02eb]=16'hffff;
      mem1[16'h02eb]=16'hffff;
      mem0[16'h02ec]=16'hffff;
      mem1[16'h02ec]=16'hffff;
      mem0[16'h02ed]=16'hffff;
      mem1[16'h02ed]=16'hffff;
      mem0[16'h02ee]=16'hffff;
      mem1[16'h02ee]=16'hffff;
      mem0[16'h02ef]=16'hffff;
      mem1[16'h02ef]=16'hffff;
      mem0[16'h02f0]=16'hffff;
      mem1[16'h02f0]=16'hffff;
      mem0[16'h02f1]=16'hffff;
      mem1[16'h02f1]=16'hffff;
      mem0[16'h02f2]=16'hffff;
      mem1[16'h02f2]=16'hffff;
      mem0[16'h02f3]=16'hffff;
      mem1[16'h02f3]=16'hffff;
      mem0[16'h02f4]=16'hffff;
      mem1[16'h02f4]=16'hffff;
      mem0[16'h02f5]=16'hffff;
      mem1[16'h02f5]=16'hffff;
      mem0[16'h02f6]=16'hffff;
      mem1[16'h02f6]=16'hffff;
      mem0[16'h02f7]=16'hffff;
      mem1[16'h02f7]=16'hffff;
      mem0[16'h02f8]=16'hffff;
      mem1[16'h02f8]=16'hffff;
      mem0[16'h02f9]=16'hffff;
      mem1[16'h02f9]=16'hffff;
      mem0[16'h02fa]=16'hffff;
      mem1[16'h02fa]=16'hffff;
      mem0[16'h02fb]=16'hffff;
      mem1[16'h02fb]=16'hffff;
      mem0[16'h02fc]=16'hffff;
      mem1[16'h02fc]=16'hffff;
      mem0[16'h02fd]=16'hffff;
      mem1[16'h02fd]=16'hffff;
      mem0[16'h02fe]=16'hffff;
      mem1[16'h02fe]=16'hffff;
      mem0[16'h02ff]=16'hffff;
      mem1[16'h02ff]=16'hffff;
      mem0[16'h0300]=16'hffff;
      mem1[16'h0300]=16'hffff;
      mem0[16'h0301]=16'hffff;
      mem1[16'h0301]=16'hffff;
      mem0[16'h0302]=16'hffff;
      mem1[16'h0302]=16'hffff;
      mem0[16'h0303]=16'hffff;
      mem1[16'h0303]=16'hffff;
      mem0[16'h0304]=16'hffff;
      mem1[16'h0304]=16'hffff;
      mem0[16'h0305]=16'hffff;
      mem1[16'h0305]=16'hffff;
      mem0[16'h0306]=16'hffff;
      mem1[16'h0306]=16'hffff;
      mem0[16'h0307]=16'hffff;
      mem1[16'h0307]=16'hffff;
      mem0[16'h0308]=16'hffff;
      mem1[16'h0308]=16'hffff;
      mem0[16'h0309]=16'hffff;
      mem1[16'h0309]=16'hffff;
      mem0[16'h030a]=16'hffff;
      mem1[16'h030a]=16'hffff;
      mem0[16'h030b]=16'hffff;
      mem1[16'h030b]=16'hffff;
      mem0[16'h030c]=16'hffff;
      mem1[16'h030c]=16'hffff;
      mem0[16'h030d]=16'hffff;
      mem1[16'h030d]=16'hffff;
      mem0[16'h030e]=16'hffff;
      mem1[16'h030e]=16'hffff;
      mem0[16'h030f]=16'hffff;
      mem1[16'h030f]=16'hffff;
      mem0[16'h0310]=16'hffff;
      mem1[16'h0310]=16'hffff;
      mem0[16'h0311]=16'hffff;
      mem1[16'h0311]=16'hffff;
      mem0[16'h0312]=16'hffff;
      mem1[16'h0312]=16'hffff;
      mem0[16'h0313]=16'hffff;
      mem1[16'h0313]=16'hffff;
      mem0[16'h0314]=16'hffff;
      mem1[16'h0314]=16'hffff;
      mem0[16'h0315]=16'hffff;
      mem1[16'h0315]=16'hffff;
      mem0[16'h0316]=16'hffff;
      mem1[16'h0316]=16'hffff;
      mem0[16'h0317]=16'hffff;
      mem1[16'h0317]=16'hffff;
      mem0[16'h0318]=16'hffff;
      mem1[16'h0318]=16'hffff;
      mem0[16'h0319]=16'hffff;
      mem1[16'h0319]=16'hffff;
      mem0[16'h031a]=16'hffff;
      mem1[16'h031a]=16'hffff;
      mem0[16'h031b]=16'hffff;
      mem1[16'h031b]=16'hffff;
      mem0[16'h031c]=16'hffff;
      mem1[16'h031c]=16'hffff;
      mem0[16'h031d]=16'hffff;
      mem1[16'h031d]=16'hffff;
      mem0[16'h031e]=16'hffff;
      mem1[16'h031e]=16'hffff;
      mem0[16'h031f]=16'hffff;
      mem1[16'h031f]=16'hffff;
      mem0[16'h0320]=16'hffff;
      mem1[16'h0320]=16'hffff;
      mem0[16'h0321]=16'hffff;
      mem1[16'h0321]=16'hffff;
      mem0[16'h0322]=16'hffff;
      mem1[16'h0322]=16'hffff;
      mem0[16'h0323]=16'hffff;
      mem1[16'h0323]=16'hffff;
      mem0[16'h0324]=16'hffff;
      mem1[16'h0324]=16'hffff;
      mem0[16'h0325]=16'hffff;
      mem1[16'h0325]=16'hffff;
      mem0[16'h0326]=16'hffff;
      mem1[16'h0326]=16'hffff;
      mem0[16'h0327]=16'hffff;
      mem1[16'h0327]=16'hffff;
      mem0[16'h0328]=16'hffff;
      mem1[16'h0328]=16'hffff;
      mem0[16'h0329]=16'hffff;
      mem1[16'h0329]=16'hffff;
      mem0[16'h032a]=16'hffff;
      mem1[16'h032a]=16'hffff;
      mem0[16'h032b]=16'hffff;
      mem1[16'h032b]=16'hffff;
      mem0[16'h032c]=16'hffff;
      mem1[16'h032c]=16'hffff;
      mem0[16'h032d]=16'hffff;
      mem1[16'h032d]=16'hffff;
      mem0[16'h032e]=16'hffff;
      mem1[16'h032e]=16'hffff;
      mem0[16'h032f]=16'hffff;
      mem1[16'h032f]=16'hffff;
      mem0[16'h0330]=16'hffff;
      mem1[16'h0330]=16'hffff;
      mem0[16'h0331]=16'hffff;
      mem1[16'h0331]=16'hffff;
      mem0[16'h0332]=16'hffff;
      mem1[16'h0332]=16'hffff;
      mem0[16'h0333]=16'hffff;
      mem1[16'h0333]=16'hffff;
      mem0[16'h0334]=16'hffff;
      mem1[16'h0334]=16'hffff;
      mem0[16'h0335]=16'hffff;
      mem1[16'h0335]=16'hffff;
      mem0[16'h0336]=16'hffff;
      mem1[16'h0336]=16'hffff;
      mem0[16'h0337]=16'hffff;
      mem1[16'h0337]=16'hffff;
      mem0[16'h0338]=16'hffff;
      mem1[16'h0338]=16'hffff;
      mem0[16'h0339]=16'hffff;
      mem1[16'h0339]=16'hffff;
      mem0[16'h033a]=16'hffff;
      mem1[16'h033a]=16'hffff;
      mem0[16'h033b]=16'hffff;
      mem1[16'h033b]=16'hffff;
      mem0[16'h033c]=16'hffff;
      mem1[16'h033c]=16'hffff;
      mem0[16'h033d]=16'hffff;
      mem1[16'h033d]=16'hffff;
      mem0[16'h033e]=16'hffff;
      mem1[16'h033e]=16'hffff;
      mem0[16'h033f]=16'hffff;
      mem1[16'h033f]=16'hffff;
      mem0[16'h0340]=16'hffff;
      mem1[16'h0340]=16'hffff;
      mem0[16'h0341]=16'hffff;
      mem1[16'h0341]=16'hffff;
      mem0[16'h0342]=16'hffff;
      mem1[16'h0342]=16'hffff;
      mem0[16'h0343]=16'hffff;
      mem1[16'h0343]=16'hffff;
      mem0[16'h0344]=16'hffff;
      mem1[16'h0344]=16'hffff;
      mem0[16'h0345]=16'hffff;
      mem1[16'h0345]=16'hffff;
      mem0[16'h0346]=16'hffff;
      mem1[16'h0346]=16'hffff;
      mem0[16'h0347]=16'hffff;
      mem1[16'h0347]=16'hffff;
      mem0[16'h0348]=16'hffff;
      mem1[16'h0348]=16'hffff;
      mem0[16'h0349]=16'hffff;
      mem1[16'h0349]=16'hffff;
      mem0[16'h034a]=16'hffff;
      mem1[16'h034a]=16'hffff;
      mem0[16'h034b]=16'hffff;
      mem1[16'h034b]=16'hffff;
      mem0[16'h034c]=16'hffff;
      mem1[16'h034c]=16'hffff;
      mem0[16'h034d]=16'hffff;
      mem1[16'h034d]=16'hffff;
      mem0[16'h034e]=16'hffff;
      mem1[16'h034e]=16'hffff;
      mem0[16'h034f]=16'hffff;
      mem1[16'h034f]=16'hffff;
      mem0[16'h0350]=16'hffff;
      mem1[16'h0350]=16'hffff;
      mem0[16'h0351]=16'hffff;
      mem1[16'h0351]=16'hffff;
      mem0[16'h0352]=16'hffff;
      mem1[16'h0352]=16'hffff;
      mem0[16'h0353]=16'hffff;
      mem1[16'h0353]=16'hffff;
      mem0[16'h0354]=16'hffff;
      mem1[16'h0354]=16'hffff;
      mem0[16'h0355]=16'hffff;
      mem1[16'h0355]=16'hffff;
      mem0[16'h0356]=16'hffff;
      mem1[16'h0356]=16'hffff;
      mem0[16'h0357]=16'hffff;
      mem1[16'h0357]=16'hffff;
      mem0[16'h0358]=16'hffff;
      mem1[16'h0358]=16'hffff;
      mem0[16'h0359]=16'hffff;
      mem1[16'h0359]=16'hffff;
      mem0[16'h035a]=16'hffff;
      mem1[16'h035a]=16'hffff;
      mem0[16'h035b]=16'hffff;
      mem1[16'h035b]=16'hffff;
      mem0[16'h035c]=16'hffff;
      mem1[16'h035c]=16'hffff;
      mem0[16'h035d]=16'hffff;
      mem1[16'h035d]=16'hffff;
      mem0[16'h035e]=16'hffff;
      mem1[16'h035e]=16'hffff;
      mem0[16'h035f]=16'hffff;
      mem1[16'h035f]=16'hffff;
      mem0[16'h0360]=16'hffff;
      mem1[16'h0360]=16'hffff;
      mem0[16'h0361]=16'hffff;
      mem1[16'h0361]=16'hffff;
      mem0[16'h0362]=16'hffff;
      mem1[16'h0362]=16'hffff;
      mem0[16'h0363]=16'hffff;
      mem1[16'h0363]=16'hffff;
      mem0[16'h0364]=16'hffff;
      mem1[16'h0364]=16'hffff;
      mem0[16'h0365]=16'hffff;
      mem1[16'h0365]=16'hffff;
      mem0[16'h0366]=16'hffff;
      mem1[16'h0366]=16'hffff;
      mem0[16'h0367]=16'hffff;
      mem1[16'h0367]=16'hffff;
      mem0[16'h0368]=16'hffff;
      mem1[16'h0368]=16'hffff;
      mem0[16'h0369]=16'hffff;
      mem1[16'h0369]=16'hffff;
      mem0[16'h036a]=16'hffff;
      mem1[16'h036a]=16'hffff;
      mem0[16'h036b]=16'hffff;
      mem1[16'h036b]=16'hffff;
      mem0[16'h036c]=16'hffff;
      mem1[16'h036c]=16'hffff;
      mem0[16'h036d]=16'hffff;
      mem1[16'h036d]=16'hffff;
      mem0[16'h036e]=16'hffff;
      mem1[16'h036e]=16'hffff;
      mem0[16'h036f]=16'hffff;
      mem1[16'h036f]=16'hffff;
      mem0[16'h0370]=16'hffff;
      mem1[16'h0370]=16'hffff;
      mem0[16'h0371]=16'hffff;
      mem1[16'h0371]=16'hffff;
      mem0[16'h0372]=16'hffff;
      mem1[16'h0372]=16'hffff;
      mem0[16'h0373]=16'hffff;
      mem1[16'h0373]=16'hffff;
      mem0[16'h0374]=16'hffff;
      mem1[16'h0374]=16'hffff;
      mem0[16'h0375]=16'hffff;
      mem1[16'h0375]=16'hffff;
      mem0[16'h0376]=16'hffff;
      mem1[16'h0376]=16'hffff;
      mem0[16'h0377]=16'hffff;
      mem1[16'h0377]=16'hffff;
      mem0[16'h0378]=16'hffff;
      mem1[16'h0378]=16'hffff;
      mem0[16'h0379]=16'hffff;
      mem1[16'h0379]=16'hffff;
      mem0[16'h037a]=16'hffff;
      mem1[16'h037a]=16'hffff;
      mem0[16'h037b]=16'hffff;
      mem1[16'h037b]=16'hffff;
      mem0[16'h037c]=16'hffff;
      mem1[16'h037c]=16'hffff;
      mem0[16'h037d]=16'hffff;
      mem1[16'h037d]=16'hffff;
      mem0[16'h037e]=16'hffff;
      mem1[16'h037e]=16'hffff;
      mem0[16'h037f]=16'hffff;
      mem1[16'h037f]=16'hffff;
      mem0[16'h0380]=16'hffff;
      mem1[16'h0380]=16'hffff;
      mem0[16'h0381]=16'hffff;
      mem1[16'h0381]=16'hffff;
      mem0[16'h0382]=16'hffff;
      mem1[16'h0382]=16'hffff;
      mem0[16'h0383]=16'hffff;
      mem1[16'h0383]=16'hffff;
      mem0[16'h0384]=16'hffff;
      mem1[16'h0384]=16'hffff;
      mem0[16'h0385]=16'hffff;
      mem1[16'h0385]=16'hffff;
      mem0[16'h0386]=16'hffff;
      mem1[16'h0386]=16'hffff;
      mem0[16'h0387]=16'hffff;
      mem1[16'h0387]=16'hffff;
      mem0[16'h0388]=16'hffff;
      mem1[16'h0388]=16'hffff;
      mem0[16'h0389]=16'hffff;
      mem1[16'h0389]=16'hffff;
      mem0[16'h038a]=16'hffff;
      mem1[16'h038a]=16'hffff;
      mem0[16'h038b]=16'hffff;
      mem1[16'h038b]=16'hffff;
      mem0[16'h038c]=16'hffff;
      mem1[16'h038c]=16'hffff;
      mem0[16'h038d]=16'hffff;
      mem1[16'h038d]=16'hffff;
      mem0[16'h038e]=16'hffff;
      mem1[16'h038e]=16'hffff;
      mem0[16'h038f]=16'hffff;
      mem1[16'h038f]=16'hffff;
      mem0[16'h0390]=16'hffff;
      mem1[16'h0390]=16'hffff;
      mem0[16'h0391]=16'hffff;
      mem1[16'h0391]=16'hffff;
      mem0[16'h0392]=16'hffff;
      mem1[16'h0392]=16'hffff;
      mem0[16'h0393]=16'hffff;
      mem1[16'h0393]=16'hffff;
      mem0[16'h0394]=16'hffff;
      mem1[16'h0394]=16'hffff;
      mem0[16'h0395]=16'hffff;
      mem1[16'h0395]=16'hffff;
      mem0[16'h0396]=16'hffff;
      mem1[16'h0396]=16'hffff;
      mem0[16'h0397]=16'hffff;
      mem1[16'h0397]=16'hffff;
      mem0[16'h0398]=16'hffff;
      mem1[16'h0398]=16'hffff;
      mem0[16'h0399]=16'hffff;
      mem1[16'h0399]=16'hffff;
      mem0[16'h039a]=16'hffff;
      mem1[16'h039a]=16'hffff;
      mem0[16'h039b]=16'hffff;
      mem1[16'h039b]=16'hffff;
      mem0[16'h039c]=16'hffff;
      mem1[16'h039c]=16'hffff;
      mem0[16'h039d]=16'hffff;
      mem1[16'h039d]=16'hffff;
      mem0[16'h039e]=16'hffff;
      mem1[16'h039e]=16'hffff;
      mem0[16'h039f]=16'hffff;
      mem1[16'h039f]=16'hffff;
      mem0[16'h03a0]=16'hffff;
      mem1[16'h03a0]=16'hffff;
      mem0[16'h03a1]=16'hffff;
      mem1[16'h03a1]=16'hffff;
      mem0[16'h03a2]=16'hffff;
      mem1[16'h03a2]=16'hffff;
      mem0[16'h03a3]=16'hffff;
      mem1[16'h03a3]=16'hffff;
      mem0[16'h03a4]=16'hffff;
      mem1[16'h03a4]=16'hffff;
      mem0[16'h03a5]=16'hffff;
      mem1[16'h03a5]=16'hffff;
      mem0[16'h03a6]=16'hffff;
      mem1[16'h03a6]=16'hffff;
      mem0[16'h03a7]=16'hffff;
      mem1[16'h03a7]=16'hffff;
      mem0[16'h03a8]=16'hffff;
      mem1[16'h03a8]=16'hffff;
      mem0[16'h03a9]=16'hffff;
      mem1[16'h03a9]=16'hffff;
      mem0[16'h03aa]=16'hffff;
      mem1[16'h03aa]=16'hffff;
      mem0[16'h03ab]=16'hffff;
      mem1[16'h03ab]=16'hffff;
      mem0[16'h03ac]=16'hffff;
      mem1[16'h03ac]=16'hffff;
      mem0[16'h03ad]=16'hffff;
      mem1[16'h03ad]=16'hffff;
      mem0[16'h03ae]=16'hffff;
      mem1[16'h03ae]=16'hffff;
      mem0[16'h03af]=16'hffff;
      mem1[16'h03af]=16'hffff;
      mem0[16'h03b0]=16'hffff;
      mem1[16'h03b0]=16'hffff;
      mem0[16'h03b1]=16'hffff;
      mem1[16'h03b1]=16'hffff;
      mem0[16'h03b2]=16'hffff;
      mem1[16'h03b2]=16'hffff;
      mem0[16'h03b3]=16'hffff;
      mem1[16'h03b3]=16'hffff;
      mem0[16'h03b4]=16'hffff;
      mem1[16'h03b4]=16'hffff;
      mem0[16'h03b5]=16'hffff;
      mem1[16'h03b5]=16'hffff;
      mem0[16'h03b6]=16'hffff;
      mem1[16'h03b6]=16'hffff;
      mem0[16'h03b7]=16'hffff;
      mem1[16'h03b7]=16'hffff;
      mem0[16'h03b8]=16'hffff;
      mem1[16'h03b8]=16'hffff;
      mem0[16'h03b9]=16'hffff;
      mem1[16'h03b9]=16'hffff;
      mem0[16'h03ba]=16'hffff;
      mem1[16'h03ba]=16'hffff;
      mem0[16'h03bb]=16'hffff;
      mem1[16'h03bb]=16'hffff;
      mem0[16'h03bc]=16'hffff;
      mem1[16'h03bc]=16'hffff;
      mem0[16'h03bd]=16'hffff;
      mem1[16'h03bd]=16'hffff;
      mem0[16'h03be]=16'hffff;
      mem1[16'h03be]=16'hffff;
      mem0[16'h03bf]=16'hffff;
      mem1[16'h03bf]=16'hffff;
      mem0[16'h03c0]=16'hffff;
      mem1[16'h03c0]=16'hffff;
      mem0[16'h03c1]=16'hffff;
      mem1[16'h03c1]=16'hffff;
      mem0[16'h03c2]=16'hffff;
      mem1[16'h03c2]=16'hffff;
      mem0[16'h03c3]=16'hffff;
      mem1[16'h03c3]=16'hffff;
      mem0[16'h03c4]=16'hffff;
      mem1[16'h03c4]=16'hffff;
      mem0[16'h03c5]=16'hffff;
      mem1[16'h03c5]=16'hffff;
      mem0[16'h03c6]=16'hffff;
      mem1[16'h03c6]=16'hffff;
      mem0[16'h03c7]=16'hffff;
      mem1[16'h03c7]=16'hffff;
      mem0[16'h03c8]=16'hffff;
      mem1[16'h03c8]=16'hffff;
      mem0[16'h03c9]=16'hffff;
      mem1[16'h03c9]=16'hffff;
      mem0[16'h03ca]=16'hffff;
      mem1[16'h03ca]=16'hffff;
      mem0[16'h03cb]=16'hffff;
      mem1[16'h03cb]=16'hffff;
      mem0[16'h03cc]=16'hffff;
      mem1[16'h03cc]=16'hffff;
      mem0[16'h03cd]=16'hffff;
      mem1[16'h03cd]=16'hffff;
      mem0[16'h03ce]=16'hffff;
      mem1[16'h03ce]=16'hffff;
      mem0[16'h03cf]=16'hffff;
      mem1[16'h03cf]=16'hffff;
      mem0[16'h03d0]=16'hffff;
      mem1[16'h03d0]=16'hffff;
      mem0[16'h03d1]=16'hffff;
      mem1[16'h03d1]=16'hffff;
      mem0[16'h03d2]=16'hffff;
      mem1[16'h03d2]=16'hffff;
      mem0[16'h03d3]=16'hffff;
      mem1[16'h03d3]=16'hffff;
      mem0[16'h03d4]=16'hffff;
      mem1[16'h03d4]=16'hffff;
      mem0[16'h03d5]=16'hffff;
      mem1[16'h03d5]=16'hffff;
      mem0[16'h03d6]=16'hffff;
      mem1[16'h03d6]=16'hffff;
      mem0[16'h03d7]=16'hffff;
      mem1[16'h03d7]=16'hffff;
      mem0[16'h03d8]=16'hffff;
      mem1[16'h03d8]=16'hffff;
      mem0[16'h03d9]=16'hffff;
      mem1[16'h03d9]=16'hffff;
      mem0[16'h03da]=16'hffff;
      mem1[16'h03da]=16'hffff;
      mem0[16'h03db]=16'hffff;
      mem1[16'h03db]=16'hffff;
      mem0[16'h03dc]=16'hffff;
      mem1[16'h03dc]=16'hffff;
      mem0[16'h03dd]=16'hffff;
      mem1[16'h03dd]=16'hffff;
      mem0[16'h03de]=16'hffff;
      mem1[16'h03de]=16'hffff;
      mem0[16'h03df]=16'hffff;
      mem1[16'h03df]=16'hffff;
      mem0[16'h03e0]=16'hffff;
      mem1[16'h03e0]=16'hffff;
      mem0[16'h03e1]=16'hffff;
      mem1[16'h03e1]=16'hffff;
      mem0[16'h03e2]=16'hffff;
      mem1[16'h03e2]=16'hffff;
      mem0[16'h03e3]=16'hffff;
      mem1[16'h03e3]=16'hffff;
      mem0[16'h03e4]=16'hffff;
      mem1[16'h03e4]=16'hffff;
      mem0[16'h03e5]=16'hffff;
      mem1[16'h03e5]=16'hffff;
      mem0[16'h03e6]=16'hffff;
      mem1[16'h03e6]=16'hffff;
      mem0[16'h03e7]=16'hffff;
      mem1[16'h03e7]=16'hffff;
      mem0[16'h03e8]=16'hffff;
      mem1[16'h03e8]=16'hffff;
      mem0[16'h03e9]=16'hffff;
      mem1[16'h03e9]=16'hffff;
      mem0[16'h03ea]=16'hffff;
      mem1[16'h03ea]=16'hffff;
      mem0[16'h03eb]=16'hffff;
      mem1[16'h03eb]=16'hffff;
      mem0[16'h03ec]=16'hffff;
      mem1[16'h03ec]=16'hffff;
      mem0[16'h03ed]=16'hffff;
      mem1[16'h03ed]=16'hffff;
      mem0[16'h03ee]=16'hffff;
      mem1[16'h03ee]=16'hffff;
      mem0[16'h03ef]=16'hffff;
      mem1[16'h03ef]=16'hffff;
      mem0[16'h03f0]=16'hffff;
      mem1[16'h03f0]=16'hffff;
      mem0[16'h03f1]=16'hffff;
      mem1[16'h03f1]=16'hffff;
      mem0[16'h03f2]=16'hffff;
      mem1[16'h03f2]=16'hffff;
      mem0[16'h03f3]=16'hffff;
      mem1[16'h03f3]=16'hffff;
      mem0[16'h03f4]=16'hffff;
      mem1[16'h03f4]=16'hffff;
      mem0[16'h03f5]=16'hffff;
      mem1[16'h03f5]=16'hffff;
      mem0[16'h03f6]=16'hffff;
      mem1[16'h03f6]=16'hffff;
      mem0[16'h03f7]=16'hffff;
      mem1[16'h03f7]=16'hffff;
      mem0[16'h03f8]=16'hffff;
      mem1[16'h03f8]=16'hffff;
      mem0[16'h03f9]=16'hffff;
      mem1[16'h03f9]=16'hffff;
      mem0[16'h03fa]=16'hffff;
      mem1[16'h03fa]=16'hffff;
      mem0[16'h03fb]=16'hffff;
      mem1[16'h03fb]=16'hffff;
      mem0[16'h03fc]=16'hffff;
      mem1[16'h03fc]=16'hffff;
      mem0[16'h03fd]=16'hffff;
      mem1[16'h03fd]=16'hffff;
      mem0[16'h03fe]=16'hffff;
      mem1[16'h03fe]=16'hffff;
      mem0[16'h03ff]=16'hffff;
      mem1[16'h03ff]=16'hffff;
      mem0[16'h0400]=16'h0000;
end
