   `include "h80cpu.svh"
   `include "h80cpu_instmacros.svh"
   initial begin
      mem[16'h0000]=16'h0160;
      mem[16'h0001]=16'h0100;
      mem[16'h0002]=16'h01e0;
      mem[16'h0003]=16'hffff;
      mem[16'h0004]=16'hffff;
      mem[16'h0005]=16'hffff;
      mem[16'h0006]=16'hffff;
      mem[16'h0007]=16'hffff;
      mem[16'h0008]=16'h0160;
      mem[16'h0009]=16'h0ab6;
      mem[16'h000a]=16'h01e0;
      mem[16'h000b]=16'hffff;
      mem[16'h000c]=16'h0160;
      mem[16'h000d]=16'h0ad2;
      mem[16'h000e]=16'h01e0;
      mem[16'h000f]=16'hffff;
      mem[16'h0010]=16'hffff;
      mem[16'h0011]=16'hffff;
      mem[16'h0012]=16'hffff;
      mem[16'h0013]=16'hffff;
      mem[16'h0014]=16'hffff;
      mem[16'h0015]=16'hffff;
      mem[16'h0016]=16'hffff;
      mem[16'h0017]=16'hffff;
      mem[16'h0018]=16'h0160;
      mem[16'h0019]=16'h0a30;
      mem[16'h001a]=16'h01e0;
      mem[16'h001b]=16'hffff;
      mem[16'h001c]=16'h0160;
      mem[16'h001d]=16'h0a32;
      mem[16'h001e]=16'h01e0;
      mem[16'h001f]=16'hffff;
      mem[16'h0020]=16'hffff;
      mem[16'h0021]=16'hffff;
      mem[16'h0022]=16'hffff;
      mem[16'h0023]=16'hffff;
      mem[16'h0024]=16'hffff;
      mem[16'h0025]=16'hffff;
      mem[16'h0026]=16'hffff;
      mem[16'h0027]=16'hffff;
      mem[16'h0028]=16'hffff;
      mem[16'h0029]=16'hffff;
      mem[16'h002a]=16'hffff;
      mem[16'h002b]=16'hffff;
      mem[16'h002c]=16'hffff;
      mem[16'h002d]=16'hffff;
      mem[16'h002e]=16'hffff;
      mem[16'h002f]=16'hffff;
      mem[16'h0030]=16'hffff;
      mem[16'h0031]=16'hffff;
      mem[16'h0032]=16'hffff;
      mem[16'h0033]=16'hffff;
      mem[16'h0034]=16'hffff;
      mem[16'h0035]=16'hffff;
      mem[16'h0036]=16'hffff;
      mem[16'h0037]=16'hffff;
      mem[16'h0038]=16'hffff;
      mem[16'h0039]=16'hffff;
      mem[16'h003a]=16'hffff;
      mem[16'h003b]=16'hffff;
      mem[16'h003c]=16'hffff;
      mem[16'h003d]=16'hffff;
      mem[16'h003e]=16'hffff;
      mem[16'h003f]=16'hffff;
      mem[16'h0040]=16'h0160;
      mem[16'h0041]=16'h0100;
      mem[16'h0042]=16'h01e0;
      mem[16'h0043]=16'hffff;
      mem[16'h0044]=16'h0160;
      mem[16'h0045]=16'h01fa;
      mem[16'h0046]=16'h01e0;
      mem[16'h0047]=16'hffff;
      mem[16'h0048]=16'h0160;
      mem[16'h0049]=16'h0ad2;
      mem[16'h004a]=16'h01e0;
      mem[16'h004b]=16'hffff;
      mem[16'h004c]=16'h0160;
      mem[16'h004d]=16'h087a;
      mem[16'h004e]=16'h01e0;
      mem[16'h004f]=16'hffff;
      mem[16'h0050]=16'h0160;
      mem[16'h0051]=16'h0ab6;
      mem[16'h0052]=16'h01e0;
      mem[16'h0053]=16'hffff;
      mem[16'h0054]=16'h0160;
      mem[16'h0055]=16'h0ac8;
      mem[16'h0056]=16'h01e0;
      mem[16'h0057]=16'hffff;
      mem[16'h0058]=16'hffff;
      mem[16'h0059]=16'hffff;
      mem[16'h005a]=16'hffff;
      mem[16'h005b]=16'hffff;
      mem[16'h005c]=16'hffff;
      mem[16'h005d]=16'hffff;
      mem[16'h005e]=16'hffff;
      mem[16'h005f]=16'hffff;
      mem[16'h0060]=16'hffff;
      mem[16'h0061]=16'hffff;
      mem[16'h0062]=16'hffff;
      mem[16'h0063]=16'hffff;
      mem[16'h0064]=16'hffff;
      mem[16'h0065]=16'hffff;
      mem[16'h0066]=16'hffff;
      mem[16'h0067]=16'hffff;
      mem[16'h0068]=16'hffff;
      mem[16'h0069]=16'hffff;
      mem[16'h006a]=16'hffff;
      mem[16'h006b]=16'hffff;
      mem[16'h006c]=16'hffff;
      mem[16'h006d]=16'hffff;
      mem[16'h006e]=16'hffff;
      mem[16'h006f]=16'hffff;
      mem[16'h0070]=16'hffff;
      mem[16'h0071]=16'hffff;
      mem[16'h0072]=16'hffff;
      mem[16'h0073]=16'hffff;
      mem[16'h0074]=16'hffff;
      mem[16'h0075]=16'hffff;
      mem[16'h0076]=16'hffff;
      mem[16'h0077]=16'hffff;
      mem[16'h0078]=16'hffff;
      mem[16'h0079]=16'hffff;
      mem[16'h007a]=16'hffff;
      mem[16'h007b]=16'hffff;
      mem[16'h007c]=16'hffff;
      mem[16'h007d]=16'hffff;
      mem[16'h007e]=16'hffff;
      mem[16'h007f]=16'hffff;
      mem[16'h0080]=16'h0166;
      mem[16'h0081]=16'h0ff0;
      mem[16'h0082]=16'h3f26;
      mem[16'h0083]=16'h0169;
      mem[16'h0084]=16'h1000;
      mem[16'h0085]=16'h016a;
      mem[16'h0086]=16'h1001;
      mem[16'h0087]=16'he666;
      mem[16'h0088]=16'he777;
      mem[16'h0089]=16'h3a6a;
      mem[16'h008a]=16'h3c67;
      mem[16'h008b]=16'h0146;
      mem[16'h008c]=16'h10ff;
      mem[16'h008d]=16'hc660;
      mem[16'h008e]=16'h386a;
      mem[16'h008f]=16'h3a4a;
      mem[16'h0090]=16'hf664;
      mem[16'h0091]=16'h0170;
      mem[16'h0092]=16'h001a;
      mem[16'h0093]=16'h0380;
      mem[16'h0094]=16'h3269;
      mem[16'h0095]=16'hf664;
      mem[16'h0096]=16'h0170;
      mem[16'h0097]=16'h001c;
      mem[16'h0098]=16'h0380;
      mem[16'h0099]=16'h307a;
      mem[16'h009a]=16'h3269;
      mem[16'h009b]=16'h3a4a;
      mem[16'h009c]=16'hf664;
      mem[16'h009d]=16'h0170;
      mem[16'h009e]=16'h000e;
      mem[16'h009f]=16'h0380;
      mem[16'h00a0]=16'h0160;
      mem[16'h00a1]=16'h0f1e;
      mem[16'h00a2]=16'h30a0;
      mem[16'h00a3]=16'h0170;
      mem[16'h00a4]=16'h0018;
      mem[16'h00a5]=16'h01f0;
      mem[16'h00a6]=16'h307a;
      mem[16'h00a7]=16'h08a1;
      mem[16'h00a8]=16'h0160;
      mem[16'h00a9]=16'h2000;
      mem[16'h00aa]=16'hfaa0;
      mem[16'h00ab]=16'h0170;
      mem[16'h00ac]=16'hffb8;
      mem[16'h00ad]=16'h03d0;
      mem[16'h00ae]=16'h0160;
      mem[16'h00af]=16'h0f1e;
      mem[16'h00b0]=16'h34a0;
      mem[16'h00b1]=16'he666;
      mem[16'h00b2]=16'h0160;
      mem[16'h00b3]=16'h0f1b;
      mem[16'h00b4]=16'h3860;
      mem[16'h00b5]=16'h0168;
      mem[16'h00b6]=16'h0a9f;
      mem[16'h00b7]=16'he999;
      mem[16'h00b8]=16'h0160;
      mem[16'h00b9]=16'h0176;
      mem[16'h00ba]=16'h01e0;
      mem[16'h00bb]=16'h0160;
      mem[16'h00bc]=16'h0f1b;
      mem[16'h00bd]=16'h3890;
      mem[16'h00be]=16'h0160;
      mem[16'h00bf]=16'h0f00;
      mem[16'h00c0]=16'h3480;
      mem[16'h00c1]=16'h0160;
      mem[16'h00c2]=16'h0ab4;
      mem[16'h00c3]=16'h01c0;
      mem[16'h00c4]=16'h0166;
      mem[16'h00c5]=16'h1000;
      mem[16'h00c6]=16'h0160;
      mem[16'h00c7]=16'h0f10;
      mem[16'h00c8]=16'h3460;
      mem[16'h00c9]=16'h0160;
      mem[16'h00ca]=16'h0f17;
      mem[16'h00cb]=16'h3460;
      mem[16'h00cc]=16'h0160;
      mem[16'h00cd]=16'h0f15;
      mem[16'h00ce]=16'h3460;
      mem[16'h00cf]=16'h1649;
      mem[16'h00d0]=16'h0160;
      mem[16'h00d1]=16'h0f19;
      mem[16'h00d2]=16'h3860;
      mem[16'h00d3]=16'he666;
      mem[16'h00d4]=16'h0160;
      mem[16'h00d5]=16'h0f1d;
      mem[16'h00d6]=16'h3860;
      mem[16'h00d7]=16'h1864;
      mem[16'h00d8]=16'he222;
      mem[16'h00d9]=16'h0160;
      mem[16'h00da]=16'h0ad2;
      mem[16'h00db]=16'h01c0;
      mem[16'h00dc]=16'h0170;
      mem[16'h00dd]=16'hfff4;
      mem[16'h00de]=16'h0a80;
      mem[16'h00df]=16'h0164;
      mem[16'h00e0]=16'h0a34;
      mem[16'h00e1]=16'h0160;
      mem[16'h00e2]=16'h087a;
      mem[16'h00e3]=16'h01c0;
      mem[16'h00e4]=16'h0160;
      mem[16'h00e5]=16'h0f00;
      mem[16'h00e6]=16'h3640;
      mem[16'h00e7]=16'h0160;
      mem[16'h00e8]=16'h087a;
      mem[16'h00e9]=16'h01c0;
      mem[16'h00ea]=16'h0164;
      mem[16'h00eb]=16'h1000;
      mem[16'h00ec]=16'h0160;
      mem[16'h00ed]=16'h088e;
      mem[16'h00ee]=16'h01c0;
      mem[16'h00ef]=16'h122d;
      mem[16'h00f0]=16'h0160;
      mem[16'h00f1]=16'h0ad2;
      mem[16'h00f2]=16'h01c0;
      mem[16'h00f3]=16'h0160;
      mem[16'h00f4]=16'h0f1e;
      mem[16'h00f5]=16'h3640;
      mem[16'h00f6]=16'h0941;
      mem[16'h00f7]=16'h0160;
      mem[16'h00f8]=16'h088e;
      mem[16'h00f9]=16'h01c0;
      mem[16'h00fa]=16'h0160;
      mem[16'h00fb]=16'h090e;
      mem[16'h00fc]=16'h01c0;
      mem[16'h00fd]=16'h0164;
      mem[16'h00fe]=16'h0a4e;
      mem[16'h00ff]=16'h0160;
      mem[16'h0100]=16'h087a;
      mem[16'h0101]=16'h01c0;
      mem[16'h0102]=16'h0160;
      mem[16'h0103]=16'h091e;
      mem[16'h0104]=16'h01c0;
      mem[16'h0105]=16'h0164;
      mem[16'h0106]=16'h0f00;
      mem[16'h0107]=16'h0160;
      mem[16'h0108]=16'h09c0;
      mem[16'h0109]=16'h01c0;
      mem[16'h010a]=16'h0160;
      mem[16'h010b]=16'h09d2;
      mem[16'h010c]=16'h01c0;
      mem[16'h010d]=16'hd222;
      mem[16'h010e]=16'h0170;
      mem[16'h010f]=16'hffda;
      mem[16'h0110]=16'h03c0;
      mem[16'h0111]=16'h1044;
      mem[16'h0112]=16'hf220;
      mem[16'h0113]=16'h0170;
      mem[16'h0114]=16'h003a;
      mem[16'h0115]=16'h03c0;
      mem[16'h0116]=16'h1047;
      mem[16'h0117]=16'hf220;
      mem[16'h0118]=16'h0160;
      mem[16'h0119]=16'h0442;
      mem[16'h011a]=16'h0340;
      mem[16'h011b]=16'h1053;
      mem[16'h011c]=16'hf220;
      mem[16'h011d]=16'h0160;
      mem[16'h011e]=16'h0474;
      mem[16'h011f]=16'h0340;
      mem[16'h0120]=16'h104c;
      mem[16'h0121]=16'hf220;
      mem[16'h0122]=16'h0160;
      mem[16'h0123]=16'h0542;
      mem[16'h0124]=16'h0340;
      mem[16'h0125]=16'h1050;
      mem[16'h0126]=16'hf220;
      mem[16'h0127]=16'h0160;
      mem[16'h0128]=16'h06e8;
      mem[16'h0129]=16'h0340;
      mem[16'h012a]=16'h0164;
      mem[16'h012b]=16'h0a6b;
      mem[16'h012c]=16'h0160;
      mem[16'h012d]=16'h087a;
      mem[16'h012e]=16'h01c0;
      mem[16'h012f]=16'h0170;
      mem[16'h0130]=16'hff98;
      mem[16'h0131]=16'h01f0;
      mem[16'h0132]=16'h0841;
      mem[16'h0133]=16'h0160;
      mem[16'h0134]=16'h09c0;
      mem[16'h0135]=16'h01c0;
      mem[16'h0136]=16'h0160;
      mem[16'h0137]=16'h09e4;
      mem[16'h0138]=16'h01c0;
      mem[16'h0139]=16'hd333;
      mem[16'h013a]=16'h0170;
      mem[16'h013b]=16'h0026;
      mem[16'h013c]=16'h0380;
      mem[16'h013d]=16'h0160;
      mem[16'h013e]=16'h09c0;
      mem[16'h013f]=16'h01c0;
      mem[16'h0140]=16'hd222;
      mem[16'h0141]=16'h0170;
      mem[16'h0142]=16'hffce;
      mem[16'h0143]=16'h0380;
      mem[16'h0144]=16'h0160;
      mem[16'h0145]=16'h0f10;
      mem[16'h0146]=16'h3660;
      mem[16'h0147]=16'h1080;
      mem[16'h0148]=16'h8660;
      mem[16'h0149]=16'h0160;
      mem[16'h014a]=16'h0f12;
      mem[16'h014b]=16'h3460;
      mem[16'h014c]=16'h0170;
      mem[16'h014d]=16'h005c;
      mem[16'h014e]=16'h01f0;
      mem[16'h014f]=16'h0160;
      mem[16'h0150]=16'h0f10;
      mem[16'h0151]=16'h3450;
      mem[16'h0152]=16'h0160;
      mem[16'h0153]=16'h09c0;
      mem[16'h0154]=16'h01c0;
      mem[16'h0155]=16'h102c;
      mem[16'h0156]=16'hf220;
      mem[16'h0157]=16'h0170;
      mem[16'h0158]=16'h001a;
      mem[16'h0159]=16'h03c0;
      mem[16'h015a]=16'hd222;
      mem[16'h015b]=16'h0170;
      mem[16'h015c]=16'hff9a;
      mem[16'h015d]=16'h0380;
      mem[16'h015e]=16'h1080;
      mem[16'h015f]=16'h8550;
      mem[16'h0160]=16'h0160;
      mem[16'h0161]=16'h0f12;
      mem[16'h0162]=16'h3450;
      mem[16'h0163]=16'h0170;
      mem[16'h0164]=16'h002e;
      mem[16'h0165]=16'h01f0;
      mem[16'h0166]=16'h0841;
      mem[16'h0167]=16'h0160;
      mem[16'h0168]=16'h09c0;
      mem[16'h0169]=16'h01c0;
      mem[16'h016a]=16'h0160;
      mem[16'h016b]=16'h09e4;
      mem[16'h016c]=16'h01c0;
      mem[16'h016d]=16'h0160;
      mem[16'h016e]=16'h09c0;
      mem[16'h016f]=16'h01c0;
      mem[16'h0170]=16'hd333;
      mem[16'h0171]=16'h0170;
      mem[16'h0172]=16'hff6e;
      mem[16'h0173]=16'h03c0;
      mem[16'h0174]=16'hd222;
      mem[16'h0175]=16'h0160;
      mem[16'h0176]=16'h0254;
      mem[16'h0177]=16'h0300;
      mem[16'h0178]=16'h0851;
      mem[16'h0179]=16'h0160;
      mem[16'h017a]=16'h0f12;
      mem[16'h017b]=16'h3450;
      mem[16'h017c]=16'he444;
      mem[16'h017d]=16'h0160;
      mem[16'h017e]=16'h0f10;
      mem[16'h017f]=16'h3640;
      mem[16'h0180]=16'h0160;
      mem[16'h0181]=16'hfff0;
      mem[16'h0182]=16'hc440;
      mem[16'h0183]=16'he666;
      mem[16'h0184]=16'h0160;
      mem[16'h0185]=16'h0f14;
      mem[16'h0186]=16'h3860;
      mem[16'h0187]=16'h0104;
      mem[16'h0188]=16'h0160;
      mem[16'h0189]=16'h035c;
      mem[16'h018a]=16'h01c0;
      mem[16'h018b]=16'h0114;
      mem[16'h018c]=16'h1010;
      mem[16'h018d]=16'h8440;
      mem[16'h018e]=16'h0160;
      mem[16'h018f]=16'h0ac8;
      mem[16'h0190]=16'h01c0;
      mem[16'h0191]=16'h0170;
      mem[16'h0192]=16'h0024;
      mem[16'h0193]=16'h0380;
      mem[16'h0194]=16'h0160;
      mem[16'h0195]=16'h0f14;
      mem[16'h0196]=16'h3a20;
      mem[16'h0197]=16'h1002;
      mem[16'h0198]=16'hf220;
      mem[16'h0199]=16'h0170;
      mem[16'h019a]=16'hffd8;
      mem[16'h019b]=16'h03d0;
      mem[16'h019c]=16'h0160;
      mem[16'h019d]=16'h0f12;
      mem[16'h019e]=16'h3240;
      mem[16'h019f]=16'h0160;
      mem[16'h01a0]=16'h0f10;
      mem[16'h01a1]=16'h3040;
      mem[16'h01a2]=16'h0160;
      mem[16'h01a3]=16'h01fa;
      mem[16'h01a4]=16'h01e0;
      mem[16'h01a5]=16'h0160;
      mem[16'h01a6]=16'h0f10;
      mem[16'h01a7]=16'h3440;
      mem[16'h01a8]=16'h0160;
      mem[16'h01a9]=16'h0ab6;
      mem[16'h01aa]=16'h01c0;
      mem[16'h01ab]=16'h0160;
      mem[16'h01ac]=16'h01fa;
      mem[16'h01ad]=16'h01e0;
      mem[16'h01ae]=16'h0160;
      mem[16'h01af]=16'h088e;
      mem[16'h01b0]=16'h01c0;
      mem[16'h01b1]=16'h0104;
      mem[16'h01b2]=16'h0164;
      mem[16'h01b3]=16'h0a73;
      mem[16'h01b4]=16'h0160;
      mem[16'h01b5]=16'h087a;
      mem[16'h01b6]=16'h01c0;
      mem[16'h01b7]=16'h0114;
      mem[16'h01b8]=16'h0168;
      mem[16'h01b9]=16'h0f00;
      mem[16'h01ba]=16'h1910;
      mem[16'h01bb]=16'h0160;
      mem[16'h01bc]=16'h03ca;
      mem[16'h01bd]=16'h01c0;
      mem[16'h01be]=16'h0170;
      mem[16'h01bf]=16'hfff6;
      mem[16'h01c0]=16'h0a90;
      mem[16'h01c1]=16'h0164;
      mem[16'h01c2]=16'h0a76;
      mem[16'h01c3]=16'h0160;
      mem[16'h01c4]=16'h087a;
      mem[16'h01c5]=16'h01c0;
      mem[16'h01c6]=16'h0164;
      mem[16'h01c7]=16'h0f00;
      mem[16'h01c8]=16'h1910;
      mem[16'h01c9]=16'h3a24;
      mem[16'h01ca]=16'h0841;
      mem[16'h01cb]=16'h1020;
      mem[16'h01cc]=16'hf220;
      mem[16'h01cd]=16'h0170;
      mem[16'h01ce]=16'h0018;
      mem[16'h01cf]=16'h03d0;
      mem[16'h01d0]=16'h107f;
      mem[16'h01d1]=16'hf220;
      mem[16'h01d2]=16'h0170;
      mem[16'h01d3]=16'h000e;
      mem[16'h01d4]=16'h0390;
      mem[16'h01d5]=16'h0160;
      mem[16'h01d6]=16'h0ad2;
      mem[16'h01d7]=16'h01c0;
      mem[16'h01d8]=16'h0170;
      mem[16'h01d9]=16'h000a;
      mem[16'h01da]=16'h01f0;
      mem[16'h01db]=16'h122e;
      mem[16'h01dc]=16'h0160;
      mem[16'h01dd]=16'h0ad2;
      mem[16'h01de]=16'h01c0;
      mem[16'h01df]=16'h0170;
      mem[16'h01e0]=16'hffd0;
      mem[16'h01e1]=16'h0a90;
      mem[16'h01e2]=16'h0160;
      mem[16'h01e3]=16'h090e;
      mem[16'h01e4]=16'h01e0;
      mem[16'h01e5]=16'h1220;
      mem[16'h01e6]=16'h0160;
      mem[16'h01e7]=16'h0ad2;
      mem[16'h01e8]=16'h01c0;
      mem[16'h01e9]=16'he666;
      mem[16'h01ea]=16'h0160;
      mem[16'h01eb]=16'h0f14;
      mem[16'h01ec]=16'h3a60;
      mem[16'h01ed]=16'hd666;
      mem[16'h01ee]=16'h0170;
      mem[16'h01ef]=16'h0030;
      mem[16'h01f0]=16'h0380;
      mem[16'h01f1]=16'he666;
      mem[16'h01f2]=16'h0160;
      mem[16'h01f3]=16'h0f10;
      mem[16'h01f4]=16'h3660;
      mem[16'h01f5]=16'hf664;
      mem[16'h01f6]=16'h0170;
      mem[16'h01f7]=16'h0018;
      mem[16'h01f8]=16'h03c0;
      mem[16'h01f9]=16'h1220;
      mem[16'h01fa]=16'h0160;
      mem[16'h01fb]=16'h0ad2;
      mem[16'h01fc]=16'h01c0;
      mem[16'h01fd]=16'h0160;
      mem[16'h01fe]=16'h0ad2;
      mem[16'h01ff]=16'h01c0;
      mem[16'h0200]=16'h3828;
      mem[16'h0201]=16'h0841;
      mem[16'h0202]=16'h0881;
      mem[16'h0203]=16'h0002;
      mem[16'h0204]=16'h1601;
      mem[16'h0205]=16'h0160;
      mem[16'h0206]=16'h0f14;
      mem[16'h0207]=16'h3860;
      mem[16'h0208]=16'h0160;
      mem[16'h0209]=16'h0f14;
      mem[16'h020a]=16'h3a60;
      mem[16'h020b]=16'h1001;
      mem[16'h020c]=16'hf660;
      mem[16'h020d]=16'h0170;
      mem[16'h020e]=16'hffd4;
      mem[16'h020f]=16'h0380;
      mem[16'h0210]=16'h3a24;
      mem[16'h0211]=16'h3828;
      mem[16'h0212]=16'h0160;
      mem[16'h0213]=16'h089a;
      mem[16'h0214]=16'h01c0;
      mem[16'h0215]=16'h0841;
      mem[16'h0216]=16'h0881;
      mem[16'h0217]=16'h0160;
      mem[16'h0218]=16'h0f12;
      mem[16'h0219]=16'h3660;
      mem[16'h021a]=16'hf446;
      mem[16'h021b]=16'h0080;
      mem[16'h021c]=16'h1602;
      mem[16'h021d]=16'h0160;
      mem[16'h021e]=16'h0f14;
      mem[16'h021f]=16'h3860;
      mem[16'h0220]=16'h0002;
      mem[16'h0221]=16'h0841;
      mem[16'h0222]=16'h0160;
      mem[16'h0223]=16'h09c0;
      mem[16'h0224]=16'h01c0;
      mem[16'h0225]=16'h0160;
      mem[16'h0226]=16'h09e4;
      mem[16'h0227]=16'h01c0;
      mem[16'h0228]=16'h0160;
      mem[16'h0229]=16'h09c0;
      mem[16'h022a]=16'h01c0;
      mem[16'h022b]=16'hd222;
      mem[16'h022c]=16'h0160;
      mem[16'h022d]=16'h0254;
      mem[16'h022e]=16'h0300;
      mem[16'h022f]=16'hd333;
      mem[16'h0230]=16'h0170;
      mem[16'h0231]=16'h0008;
      mem[16'h0232]=16'h03c0;
      mem[16'h0233]=16'h0160;
      mem[16'h0234]=16'h0f15;
      mem[16'h0235]=16'h3450;
      mem[16'h0236]=16'h0160;
      mem[16'h0237]=16'h0f15;
      mem[16'h0238]=16'h3660;
      mem[16'h0239]=16'h01e6;
      mem[16'h023a]=16'h0841;
      mem[16'h023b]=16'h0160;
      mem[16'h023c]=16'h09c0;
      mem[16'h023d]=16'h01c0;
      mem[16'h023e]=16'h0160;
      mem[16'h023f]=16'h09e4;
      mem[16'h0240]=16'h01c0;
      mem[16'h0241]=16'h0160;
      mem[16'h0242]=16'h09c0;
      mem[16'h0243]=16'h01c0;
      mem[16'h0244]=16'hd222;
      mem[16'h0245]=16'h0160;
      mem[16'h0246]=16'h0254;
      mem[16'h0247]=16'h0300;
      mem[16'h0248]=16'hd333;
      mem[16'h0249]=16'h0170;
      mem[16'h024a]=16'h000a;
      mem[16'h024b]=16'h0380;
      mem[16'h024c]=16'he555;
      mem[16'h024d]=16'h0160;
      mem[16'h024e]=16'h0f17;
      mem[16'h024f]=16'h3650;
      mem[16'h0250]=16'h0c45;
      mem[16'h0251]=16'h0160;
      mem[16'h0252]=16'h088e;
      mem[16'h0253]=16'h01c0;
      mem[16'h0254]=16'h0104;
      mem[16'h0255]=16'h0164;
      mem[16'h0256]=16'h0a76;
      mem[16'h0257]=16'h0160;
      mem[16'h0258]=16'h087a;
      mem[16'h0259]=16'h01c0;
      mem[16'h025a]=16'h0114;
      mem[16'h025b]=16'h3a24;
      mem[16'h025c]=16'h0104;
      mem[16'h025d]=16'h0160;
      mem[16'h025e]=16'h089a;
      mem[16'h025f]=16'h01c0;
      mem[16'h0260]=16'h1220;
      mem[16'h0261]=16'h0160;
      mem[16'h0262]=16'h0ad2;
      mem[16'h0263]=16'h01c0;
      mem[16'h0264]=16'h0160;
      mem[16'h0265]=16'h091e;
      mem[16'h0266]=16'h01c0;
      mem[16'h0267]=16'h0164;
      mem[16'h0268]=16'h0f00;
      mem[16'h0269]=16'h0160;
      mem[16'h026a]=16'h09c0;
      mem[16'h026b]=16'h01c0;
      mem[16'h026c]=16'hd222;
      mem[16'h026d]=16'h0170;
      mem[16'h026e]=16'h0012;
      mem[16'h026f]=16'h0380;
      mem[16'h0270]=16'h0114;
      mem[16'h0271]=16'h0841;
      mem[16'h0272]=16'h0160;
      mem[16'h0273]=16'h0f17;
      mem[16'h0274]=16'h3040;
      mem[16'h0275]=16'h0170;
      mem[16'h0276]=16'hffb4;
      mem[16'h0277]=16'h01f0;
      mem[16'h0278]=16'h102d;
      mem[16'h0279]=16'hf220;
      mem[16'h027a]=16'h0170;
      mem[16'h027b]=16'h0012;
      mem[16'h027c]=16'h0380;
      mem[16'h027d]=16'h0114;
      mem[16'h027e]=16'h0941;
      mem[16'h027f]=16'h0160;
      mem[16'h0280]=16'h0f17;
      mem[16'h0281]=16'h3040;
      mem[16'h0282]=16'h0170;
      mem[16'h0283]=16'hff9a;
      mem[16'h0284]=16'h01f0;
      mem[16'h0285]=16'h102e;
      mem[16'h0286]=16'hf220;
      mem[16'h0287]=16'h0170;
      mem[16'h0288]=16'h0010;
      mem[16'h0289]=16'h0380;
      mem[16'h028a]=16'h0114;
      mem[16'h028b]=16'h0160;
      mem[16'h028c]=16'h0f17;
      mem[16'h028d]=16'h3040;
      mem[16'h028e]=16'h0160;
      mem[16'h028f]=16'h01fa;
      mem[16'h0290]=16'h01e0;
      mem[16'h0291]=16'h0160;
      mem[16'h0292]=16'h09e4;
      mem[16'h0293]=16'h01c0;
      mem[16'h0294]=16'hd333;
      mem[16'h0295]=16'h0114;
      mem[16'h0296]=16'h0160;
      mem[16'h0297]=16'h0254;
      mem[16'h0298]=16'h0340;
      mem[16'h0299]=16'h3854;
      mem[16'h029a]=16'h0841;
      mem[16'h029b]=16'h0160;
      mem[16'h029c]=16'h0f17;
      mem[16'h029d]=16'h3040;
      mem[16'h029e]=16'h0170;
      mem[16'h029f]=16'hff62;
      mem[16'h02a0]=16'h01f0;
      mem[16'h02a1]=16'h0841;
      mem[16'h02a2]=16'h0160;
      mem[16'h02a3]=16'h09c0;
      mem[16'h02a4]=16'h01c0;
      mem[16'h02a5]=16'h0160;
      mem[16'h02a6]=16'h09e4;
      mem[16'h02a7]=16'h01c0;
      mem[16'h02a8]=16'h0160;
      mem[16'h02a9]=16'h09c0;
      mem[16'h02aa]=16'h01c0;
      mem[16'h02ab]=16'hd222;
      mem[16'h02ac]=16'h0160;
      mem[16'h02ad]=16'h0254;
      mem[16'h02ae]=16'h0300;
      mem[16'h02af]=16'hd333;
      mem[16'h02b0]=16'h0170;
      mem[16'h02b1]=16'h0004;
      mem[16'h02b2]=16'h0380;
      mem[16'h02b3]=16'h1500;
      mem[16'h02b4]=16'h0160;
      mem[16'h02b5]=16'h0ab6;
      mem[16'h02b6]=16'h01c0;
      mem[16'h02b7]=16'h0160;
      mem[16'h02b8]=16'h09d2;
      mem[16'h02b9]=16'h01c0;
      mem[16'h02ba]=16'h1053;
      mem[16'h02bb]=16'hf220;
      mem[16'h02bc]=16'h0170;
      mem[16'h02bd]=16'h00c0;
      mem[16'h02be]=16'h03c0;
      mem[16'h02bf]=16'h103a;
      mem[16'h02c0]=16'hf220;
      mem[16'h02c1]=16'h0170;
      mem[16'h02c2]=16'h0022;
      mem[16'h02c3]=16'h03c0;
      mem[16'h02c4]=16'h100d;
      mem[16'h02c5]=16'hf220;
      mem[16'h02c6]=16'h0170;
      mem[16'h02c7]=16'hffd8;
      mem[16'h02c8]=16'h03c0;
      mem[16'h02c9]=16'h100a;
      mem[16'h02ca]=16'hf220;
      mem[16'h02cb]=16'h0170;
      mem[16'h02cc]=16'hffce;
      mem[16'h02cd]=16'h03c0;
      mem[16'h02ce]=16'h0160;
      mem[16'h02cf]=16'h0ab6;
      mem[16'h02d0]=16'h01c0;
      mem[16'h02d1]=16'h0170;
      mem[16'h02d2]=16'hffe2;
      mem[16'h02d3]=16'h01f0;
      mem[16'h02d4]=16'h0160;
      mem[16'h02d5]=16'h08c0;
      mem[16'h02d6]=16'h01c0;
      mem[16'h02d7]=16'h3c29;
      mem[16'h02d8]=16'h3c28;
      mem[16'h02d9]=16'h0160;
      mem[16'h02da]=16'h08c0;
      mem[16'h02db]=16'h01c0;
      mem[16'h02dc]=16'h8992;
      mem[16'h02dd]=16'h0628;
      mem[16'h02de]=16'h3c24;
      mem[16'h02df]=16'h0160;
      mem[16'h02e0]=16'h08c0;
      mem[16'h02e1]=16'h01c0;
      mem[16'h02e2]=16'hd442;
      mem[16'h02e3]=16'h8992;
      mem[16'h02e4]=16'h8445;
      mem[16'h02e5]=16'h0160;
      mem[16'h02e6]=16'h08c0;
      mem[16'h02e7]=16'h01c0;
      mem[16'h02e8]=16'h0160;
      mem[16'h02e9]=16'h0f1a;
      mem[16'h02ea]=16'h3820;
      mem[16'h02eb]=16'h8992;
      mem[16'h02ec]=16'hd888;
      mem[16'h02ed]=16'h0170;
      mem[16'h02ee]=16'h0024;
      mem[16'h02ef]=16'h03c0;
      mem[16'h02f0]=16'h0160;
      mem[16'h02f1]=16'h08c0;
      mem[16'h02f2]=16'h01c0;
      mem[16'h02f3]=16'h8992;
      mem[16'h02f4]=16'he666;
      mem[16'h02f5]=16'h0160;
      mem[16'h02f6]=16'h0f1a;
      mem[16'h02f7]=16'h3a60;
      mem[16'h02f8]=16'hd666;
      mem[16'h02f9]=16'h0170;
      mem[16'h02fa]=16'h0006;
      mem[16'h02fb]=16'h0380;
      mem[16'h02fc]=16'h3824;
      mem[16'h02fd]=16'h0841;
      mem[16'h02fe]=16'h0170;
      mem[16'h02ff]=16'hffe0;
      mem[16'h0300]=16'h0a80;
      mem[16'h0301]=16'h0160;
      mem[16'h0302]=16'h08c0;
      mem[16'h0303]=16'h01c0;
      mem[16'h0304]=16'h8992;
      mem[16'h0305]=16'h10ff;
      mem[16'h0306]=16'hc990;
      mem[16'h0307]=16'hd999;
      mem[16'h0308]=16'h0170;
      mem[16'h0309]=16'h0018;
      mem[16'h030a]=16'h0380;
      mem[16'h030b]=16'he666;
      mem[16'h030c]=16'h0160;
      mem[16'h030d]=16'h0f1a;
      mem[16'h030e]=16'h3a60;
      mem[16'h030f]=16'hd666;
      mem[16'h0310]=16'h0160;
      mem[16'h0311]=16'h059c;
      mem[16'h0312]=16'h0340;
      mem[16'h0313]=16'h0160;
      mem[16'h0314]=16'h01fa;
      mem[16'h0315]=16'h01e0;
      mem[16'h0316]=16'h0164;
      mem[16'h0317]=16'h0a51;
      mem[16'h0318]=16'h0160;
      mem[16'h0319]=16'h087a;
      mem[16'h031a]=16'h01c0;
      mem[16'h031b]=16'h0160;
      mem[16'h031c]=16'h01fa;
      mem[16'h031d]=16'h01e0;
      mem[16'h031e]=16'h0160;
      mem[16'h031f]=16'h0ab6;
      mem[16'h0320]=16'h01c0;
      mem[16'h0321]=16'h0160;
      mem[16'h0322]=16'h0f1a;
      mem[16'h0323]=16'h3820;
      mem[16'h0324]=16'h0160;
      mem[16'h0325]=16'h08c0;
      mem[16'h0326]=16'h01c0;
      mem[16'h0327]=16'h3c28;
      mem[16'h0328]=16'h3c29;
      mem[16'h0329]=16'h0160;
      mem[16'h032a]=16'h08c0;
      mem[16'h032b]=16'h01c0;
      mem[16'h032c]=16'h8992;
      mem[16'h032d]=16'h0628;
      mem[16'h032e]=16'h3c24;
      mem[16'h032f]=16'h0160;
      mem[16'h0330]=16'h08c0;
      mem[16'h0331]=16'h01c0;
      mem[16'h0332]=16'hd442;
      mem[16'h0333]=16'h8992;
      mem[16'h0334]=16'h8445;
      mem[16'h0335]=16'h0983;
      mem[16'h0336]=16'h0170;
      mem[16'h0337]=16'h0026;
      mem[16'h0338]=16'h03c0;
      mem[16'h0339]=16'h0160;
      mem[16'h033a]=16'h08c0;
      mem[16'h033b]=16'h01c0;
      mem[16'h033c]=16'h8992;
      mem[16'h033d]=16'he666;
      mem[16'h033e]=16'h0160;
      mem[16'h033f]=16'h0f1a;
      mem[16'h0340]=16'h3a60;
      mem[16'h0341]=16'h1031;
      mem[16'h0342]=16'hf660;
      mem[16'h0343]=16'h0170;
      mem[16'h0344]=16'h0006;
      mem[16'h0345]=16'h0380;
      mem[16'h0346]=16'h3824;
      mem[16'h0347]=16'h0841;
      mem[16'h0348]=16'h0170;
      mem[16'h0349]=16'hffde;
      mem[16'h034a]=16'h0a80;
      mem[16'h034b]=16'h0160;
      mem[16'h034c]=16'h08c0;
      mem[16'h034d]=16'h01c0;
      mem[16'h034e]=16'h8992;
      mem[16'h034f]=16'h10ff;
      mem[16'h0350]=16'hc990;
      mem[16'h0351]=16'h10ff;
      mem[16'h0352]=16'hf990;
      mem[16'h0353]=16'h0170;
      mem[16'h0354]=16'h002e;
      mem[16'h0355]=16'h0380;
      mem[16'h0356]=16'he666;
      mem[16'h0357]=16'h0160;
      mem[16'h0358]=16'h0f1a;
      mem[16'h0359]=16'h3a60;
      mem[16'h035a]=16'h1037;
      mem[16'h035b]=16'hf660;
      mem[16'h035c]=16'h0170;
      mem[16'h035d]=16'h0026;
      mem[16'h035e]=16'h03c0;
      mem[16'h035f]=16'h1038;
      mem[16'h0360]=16'hf660;
      mem[16'h0361]=16'h0170;
      mem[16'h0362]=16'h001c;
      mem[16'h0363]=16'h03c0;
      mem[16'h0364]=16'h1039;
      mem[16'h0365]=16'hf660;
      mem[16'h0366]=16'h0170;
      mem[16'h0367]=16'h0012;
      mem[16'h0368]=16'h03c0;
      mem[16'h0369]=16'h0160;
      mem[16'h036a]=16'h059c;
      mem[16'h036b]=16'h01e0;
      mem[16'h036c]=16'h0164;
      mem[16'h036d]=16'h0a5e;
      mem[16'h036e]=16'h0160;
      mem[16'h036f]=16'h087a;
      mem[16'h0370]=16'h01c0;
      mem[16'h0371]=16'h0160;
      mem[16'h0372]=16'h01fa;
      mem[16'h0373]=16'h01e0;
      mem[16'h0374]=16'h0841;
      mem[16'h0375]=16'he222;
      mem[16'h0376]=16'h3a24;
      mem[16'h0377]=16'h0160;
      mem[16'h0378]=16'h09d2;
      mem[16'h0379]=16'h01c0;
      mem[16'h037a]=16'h1049;
      mem[16'h037b]=16'hf220;
      mem[16'h037c]=16'h0170;
      mem[16'h037d]=16'h000c;
      mem[16'h037e]=16'h03c0;
      mem[16'h037f]=16'h1053;
      mem[16'h0380]=16'hf220;
      mem[16'h0381]=16'h0170;
      mem[16'h0382]=16'h000a;
      mem[16'h0383]=16'h0380;
      mem[16'h0384]=16'h0841;
      mem[16'h0385]=16'h0160;
      mem[16'h0386]=16'h0f19;
      mem[16'h0387]=16'h3820;
      mem[16'h0388]=16'h0160;
      mem[16'h0389]=16'h09c0;
      mem[16'h038a]=16'h01c0;
      mem[16'h038b]=16'h0160;
      mem[16'h038c]=16'h09e4;
      mem[16'h038d]=16'h01c0;
      mem[16'h038e]=16'hd333;
      mem[16'h038f]=16'h0170;
      mem[16'h0390]=16'h0038;
      mem[16'h0391]=16'h03c0;
      mem[16'h0392]=16'h3c58;
      mem[16'h0393]=16'h0160;
      mem[16'h0394]=16'h09c0;
      mem[16'h0395]=16'h01c0;
      mem[16'h0396]=16'h102c;
      mem[16'h0397]=16'hf220;
      mem[16'h0398]=16'h0170;
      mem[16'h0399]=16'h0026;
      mem[16'h039a]=16'h0380;
      mem[16'h039b]=16'h0841;
      mem[16'h039c]=16'h0160;
      mem[16'h039d]=16'h09c0;
      mem[16'h039e]=16'h01c0;
      mem[16'h039f]=16'h0160;
      mem[16'h03a0]=16'h09e4;
      mem[16'h03a1]=16'h01c0;
      mem[16'h03a2]=16'hd333;
      mem[16'h03a3]=16'h0170;
      mem[16'h03a4]=16'h0010;
      mem[16'h03a5]=16'h03c0;
      mem[16'h03a6]=16'h0160;
      mem[16'h03a7]=16'h09c0;
      mem[16'h03a8]=16'h01c0;
      mem[16'h03a9]=16'hd222;
      mem[16'h03aa]=16'h0170;
      mem[16'h03ab]=16'h0008;
      mem[16'h03ac]=16'h03c0;
      mem[16'h03ad]=16'h0160;
      mem[16'h03ae]=16'h0254;
      mem[16'h03af]=16'h01e0;
      mem[16'h03b0]=16'h3c84;
      mem[16'h03b1]=16'h0c45;
      mem[16'h03b2]=16'h0841;
      mem[16'h03b3]=16'h9445;
      mem[16'h03b4]=16'h0160;
      mem[16'h03b5]=16'h07a8;
      mem[16'h03b6]=16'h01c0;
      mem[16'h03b7]=16'hd444;
      mem[16'h03b8]=16'h0170;
      mem[16'h03b9]=16'hfff4;
      mem[16'h03ba]=16'h0380;
      mem[16'h03bb]=16'he666;
      mem[16'h03bc]=16'h0160;
      mem[16'h03bd]=16'h0f19;
      mem[16'h03be]=16'h3a60;
      mem[16'h03bf]=16'h1049;
      mem[16'h03c0]=16'hf660;
      mem[16'h03c1]=16'h0170;
      mem[16'h03c2]=16'h0012;
      mem[16'h03c3]=16'h0380;
      mem[16'h03c4]=16'h0164;
      mem[16'h03c5]=16'h0a7a;
      mem[16'h03c6]=16'h0160;
      mem[16'h03c7]=16'h087a;
      mem[16'h03c8]=16'h01c0;
      mem[16'h03c9]=16'h0160;
      mem[16'h03ca]=16'h01fa;
      mem[16'h03cb]=16'h01e0;
      mem[16'h03cc]=16'h0164;
      mem[16'h03cd]=16'h0a88;
      mem[16'h03ce]=16'h0160;
      mem[16'h03cf]=16'h087a;
      mem[16'h03d0]=16'h01c0;
      mem[16'h03d1]=16'h0160;
      mem[16'h03d2]=16'h01fa;
      mem[16'h03d3]=16'h01e0;
      mem[16'h03d4]=16'h1810;
      mem[16'h03d5]=16'hf448;
      mem[16'h03d6]=16'h0170;
      mem[16'h03d7]=16'h0004;
      mem[16'h03d8]=16'h0390;
      mem[16'h03d9]=16'h3c48;
      mem[16'h03da]=16'h9448;
      mem[16'h03db]=16'he666;
      mem[16'h03dc]=16'h0160;
      mem[16'h03dd]=16'h0f19;
      mem[16'h03de]=16'h3a60;
      mem[16'h03df]=16'h1049;
      mem[16'h03e0]=16'hf660;
      mem[16'h03e1]=16'h0170;
      mem[16'h03e2]=16'h005a;
      mem[16'h03e3]=16'h0380;
      mem[16'h03e4]=16'h123a;
      mem[16'h03e5]=16'h0160;
      mem[16'h03e6]=16'h0ad2;
      mem[16'h03e7]=16'h01c0;
      mem[16'h03e8]=16'h3c82;
      mem[16'h03e9]=16'h0160;
      mem[16'h03ea]=16'h089a;
      mem[16'h03eb]=16'h01c0;
      mem[16'h03ec]=16'h3c89;
      mem[16'h03ed]=16'h3c52;
      mem[16'h03ee]=16'h0528;
      mem[16'h03ef]=16'h8992;
      mem[16'h03f0]=16'h0160;
      mem[16'h03f1]=16'h089a;
      mem[16'h03f2]=16'h01c0;
      mem[16'h03f3]=16'hc225;
      mem[16'h03f4]=16'h10ff;
      mem[16'h03f5]=16'hc220;
      mem[16'h03f6]=16'h8992;
      mem[16'h03f7]=16'h0160;
      mem[16'h03f8]=16'h089a;
      mem[16'h03f9]=16'h01c0;
      mem[16'h03fa]=16'he222;
      mem[16'h03fb]=16'h0160;
      mem[16'h03fc]=16'h089a;
      mem[16'h03fd]=16'h01c0;
      mem[16'h03fe]=16'he222;
      mem[16'h03ff]=16'h3a25;
      mem[16'h0400]=16'h8992;
      mem[16'h0401]=16'h0160;
      mem[16'h0402]=16'h089a;
      mem[16'h0403]=16'h01c0;
      mem[16'h0404]=16'h0851;
      mem[16'h0405]=16'h0170;
      mem[16'h0406]=16'hffee;
      mem[16'h0407]=16'h0a80;
      mem[16'h0408]=16'h0159;
      mem[16'h0409]=16'h3c92;
      mem[16'h040a]=16'h0160;
      mem[16'h040b]=16'h089a;
      mem[16'h040c]=16'h01c0;
      mem[16'h040d]=16'h0160;
      mem[16'h040e]=16'h090e;
      mem[16'h040f]=16'h01e0;
      mem[16'h0410]=16'h1253;
      mem[16'h0411]=16'h0160;
      mem[16'h0412]=16'h0ad2;
      mem[16'h0413]=16'h01c0;
      mem[16'h0414]=16'h1231;
      mem[16'h0415]=16'h0160;
      mem[16'h0416]=16'h0ad2;
      mem[16'h0417]=16'h01c0;
      mem[16'h0418]=16'h0883;
      mem[16'h0419]=16'h3c89;
      mem[16'h041a]=16'h3c82;
      mem[16'h041b]=16'h0160;
      mem[16'h041c]=16'h089a;
      mem[16'h041d]=16'h01c0;
      mem[16'h041e]=16'h3c42;
      mem[16'h041f]=16'h0528;
      mem[16'h0420]=16'h3c29;
      mem[16'h0421]=16'h0160;
      mem[16'h0422]=16'h089a;
      mem[16'h0423]=16'h01c0;
      mem[16'h0424]=16'h3c42;
      mem[16'h0425]=16'h10ff;
      mem[16'h0426]=16'hc220;
      mem[16'h0427]=16'h3c29;
      mem[16'h0428]=16'h0160;
      mem[16'h0429]=16'h089a;
      mem[16'h042a]=16'h01c0;
      mem[16'h042b]=16'he222;
      mem[16'h042c]=16'h3a25;
      mem[16'h042d]=16'h8992;
      mem[16'h042e]=16'h0160;
      mem[16'h042f]=16'h089a;
      mem[16'h0430]=16'h01c0;
      mem[16'h0431]=16'h0851;
      mem[16'h0432]=16'h0170;
      mem[16'h0433]=16'hffee;
      mem[16'h0434]=16'h0a80;
      mem[16'h0435]=16'h0149;
      mem[16'h0436]=16'h3c92;
      mem[16'h0437]=16'h0160;
      mem[16'h0438]=16'h089a;
      mem[16'h0439]=16'h01c0;
      mem[16'h043a]=16'h0160;
      mem[16'h043b]=16'h090e;
      mem[16'h043c]=16'h01e0;
      mem[16'h043d]=16'h3a24;
      mem[16'h043e]=16'hc222;
      mem[16'h043f]=16'h0084;
      mem[16'h0440]=16'h0160;
      mem[16'h0441]=16'h0ad2;
      mem[16'h0442]=16'h01c0;
      mem[16'h0443]=16'h0841;
      mem[16'h0444]=16'h0170;
      mem[16'h0445]=16'hffee;
      mem[16'h0446]=16'h01f0;
      mem[16'h0447]=16'h3c42;
      mem[16'h0448]=16'h0428;
      mem[16'h0449]=16'h0160;
      mem[16'h044a]=16'h089a;
      mem[16'h044b]=16'h01c0;
      mem[16'h044c]=16'h3c42;
      mem[16'h044d]=16'h3c26;
      mem[16'h044e]=16'h0424;
      mem[16'h044f]=16'h0160;
      mem[16'h0450]=16'h08a6;
      mem[16'h0451]=16'h01c0;
      mem[16'h0452]=16'h3c62;
      mem[16'h0453]=16'h100f;
      mem[16'h0454]=16'hc220;
      mem[16'h0455]=16'h1030;
      mem[16'h0456]=16'h8220;
      mem[16'h0457]=16'h103a;
      mem[16'h0458]=16'hf220;
      mem[16'h0459]=16'h0160;
      mem[16'h045a]=16'h0ad2;
      mem[16'h045b]=16'h0350;
      mem[16'h045c]=16'h0827;
      mem[16'h045d]=16'h0160;
      mem[16'h045e]=16'h0ad2;
      mem[16'h045f]=16'h01e0;
      mem[16'h0460]=16'he222;
      mem[16'h0461]=16'h0160;
      mem[16'h0462]=16'h08ca;
      mem[16'h0463]=16'h01c0;
      mem[16'h0464]=16'h0624;
      mem[16'h0465]=16'h0108;
      mem[16'h0466]=16'h3c28;
      mem[16'h0467]=16'h0160;
      mem[16'h0468]=16'h0ab6;
      mem[16'h0469]=16'h01c0;
      mem[16'h046a]=16'h0160;
      mem[16'h046b]=16'h09d2;
      mem[16'h046c]=16'h01c0;
      mem[16'h046d]=16'h1030;
      mem[16'h046e]=16'hf220;
      mem[16'h046f]=16'h0170;
      mem[16'h0470]=16'h0028;
      mem[16'h0471]=16'h03d0;
      mem[16'h0472]=16'h103a;
      mem[16'h0473]=16'hf220;
      mem[16'h0474]=16'h0170;
      mem[16'h0475]=16'h0018;
      mem[16'h0476]=16'h03d0;
      mem[16'h0477]=16'h1041;
      mem[16'h0478]=16'hf220;
      mem[16'h0479]=16'h0170;
      mem[16'h047a]=16'h0014;
      mem[16'h047b]=16'h03d0;
      mem[16'h047c]=16'h1047;
      mem[16'h047d]=16'hf220;
      mem[16'h047e]=16'h0170;
      mem[16'h047f]=16'h000a;
      mem[16'h0480]=16'h0390;
      mem[16'h0481]=16'h0927;
      mem[16'h0482]=16'h1030;
      mem[16'h0483]=16'h9220;
      mem[16'h0484]=16'hd228;
      mem[16'h0485]=16'h0118;
      mem[16'h0486]=16'h0002;
      mem[16'h0487]=16'h120d;
      mem[16'h0488]=16'h0160;
      mem[16'h0489]=16'h0ad2;
      mem[16'h048a]=16'h01c0;
      mem[16'h048b]=16'h120a;
      mem[16'h048c]=16'h0160;
      mem[16'h048d]=16'h0ad2;
      mem[16'h048e]=16'h01e0;
      mem[16'h048f]=16'h010a;
      mem[16'h0490]=16'h0108;
      mem[16'h0491]=16'h016a;
      mem[16'h0492]=16'h0f00;
      mem[16'h0493]=16'h1800;
      mem[16'h0494]=16'h0160;
      mem[16'h0495]=16'h0ab6;
      mem[16'h0496]=16'h01c0;
      mem[16'h0497]=16'h100d;
      mem[16'h0498]=16'hf220;
      mem[16'h0499]=16'h0170;
      mem[16'h049a]=16'h007a;
      mem[16'h049b]=16'h03c0;
      mem[16'h049c]=16'h100a;
      mem[16'h049d]=16'hf220;
      mem[16'h049e]=16'h0170;
      mem[16'h049f]=16'h0070;
      mem[16'h04a0]=16'h03c0;
      mem[16'h04a1]=16'h1008;
      mem[16'h04a2]=16'hf220;
      mem[16'h04a3]=16'h0170;
      mem[16'h04a4]=16'h003c;
      mem[16'h04a5]=16'h03c0;
      mem[16'h04a6]=16'h107f;
      mem[16'h04a7]=16'hf220;
      mem[16'h04a8]=16'h0170;
      mem[16'h04a9]=16'h0032;
      mem[16'h04aa]=16'h03c0;
      mem[16'h04ab]=16'h1020;
      mem[16'h04ac]=16'hf220;
      mem[16'h04ad]=16'h0170;
      mem[16'h04ae]=16'hffca;
      mem[16'h04af]=16'h03d0;
      mem[16'h04b0]=16'h1080;
      mem[16'h04b1]=16'hf220;
      mem[16'h04b2]=16'h0170;
      mem[16'h04b3]=16'hffc0;
      mem[16'h04b4]=16'h0390;
      mem[16'h04b5]=16'h100f;
      mem[16'h04b6]=16'hf880;
      mem[16'h04b7]=16'h0170;
      mem[16'h04b8]=16'hffb6;
      mem[16'h04b9]=16'h0390;
      mem[16'h04ba]=16'h0881;
      mem[16'h04bb]=16'h0160;
      mem[16'h04bc]=16'h0ad2;
      mem[16'h04bd]=16'h01c0;
      mem[16'h04be]=16'h382a;
      mem[16'h04bf]=16'h08a1;
      mem[16'h04c0]=16'h0170;
      mem[16'h04c1]=16'hffa4;
      mem[16'h04c2]=16'h01f0;
      mem[16'h04c3]=16'hc888;
      mem[16'h04c4]=16'h0170;
      mem[16'h04c5]=16'hff9c;
      mem[16'h04c6]=16'h03c0;
      mem[16'h04c7]=16'h0981;
      mem[16'h04c8]=16'h09a1;
      mem[16'h04c9]=16'h1208;
      mem[16'h04ca]=16'h0160;
      mem[16'h04cb]=16'h0ad2;
      mem[16'h04cc]=16'h01c0;
      mem[16'h04cd]=16'h1220;
      mem[16'h04ce]=16'h0160;
      mem[16'h04cf]=16'h0ad2;
      mem[16'h04d0]=16'h01c0;
      mem[16'h04d1]=16'h1208;
      mem[16'h04d2]=16'h0160;
      mem[16'h04d3]=16'h0ad2;
      mem[16'h04d4]=16'h01c0;
      mem[16'h04d5]=16'h0170;
      mem[16'h04d6]=16'hff7a;
      mem[16'h04d7]=16'h01f0;
      mem[16'h04d8]=16'h0160;
      mem[16'h04d9]=16'h090e;
      mem[16'h04da]=16'h01c0;
      mem[16'h04db]=16'h1000;
      mem[16'h04dc]=16'h380a;
      mem[16'h04dd]=16'h0118;
      mem[16'h04de]=16'h011a;
      mem[16'h04df]=16'h0002;
      mem[16'h04e0]=16'he222;
      mem[16'h04e1]=16'h3a24;
      mem[16'h04e2]=16'h1020;
      mem[16'h04e3]=16'hf220;
      mem[16'h04e4]=16'h0080;
      mem[16'h04e5]=16'h0841;
      mem[16'h04e6]=16'h0170;
      mem[16'h04e7]=16'hfff0;
      mem[16'h04e8]=16'h01f0;
      mem[16'h04e9]=16'h1061;
      mem[16'h04ea]=16'hf220;
      mem[16'h04eb]=16'h0085;
      mem[16'h04ec]=16'h107b;
      mem[16'h04ed]=16'hf220;
      mem[16'h04ee]=16'h0081;
      mem[16'h04ef]=16'h20e0;
      mem[16'h04f0]=16'h8220;
      mem[16'h04f1]=16'h0002;
      mem[16'h04f2]=16'he555;
      mem[16'h04f3]=16'he333;
      mem[16'h04f4]=16'he222;
      mem[16'h04f5]=16'h3a24;
      mem[16'h04f6]=16'h0160;
      mem[16'h04f7]=16'h09d2;
      mem[16'h04f8]=16'h01c0;
      mem[16'h04f9]=16'h1030;
      mem[16'h04fa]=16'hf220;
      mem[16'h04fb]=16'h0170;
      mem[16'h04fc]=16'h0034;
      mem[16'h04fd]=16'h03d0;
      mem[16'h04fe]=16'h103a;
      mem[16'h04ff]=16'hf220;
      mem[16'h0500]=16'h0170;
      mem[16'h0501]=16'h0018;
      mem[16'h0502]=16'h03d0;
      mem[16'h0503]=16'h1041;
      mem[16'h0504]=16'hf220;
      mem[16'h0505]=16'h0170;
      mem[16'h0506]=16'h0020;
      mem[16'h0507]=16'h03d0;
      mem[16'h0508]=16'h1047;
      mem[16'h0509]=16'hf220;
      mem[16'h050a]=16'h0170;
      mem[16'h050b]=16'h0016;
      mem[16'h050c]=16'h0390;
      mem[16'h050d]=16'h0927;
      mem[16'h050e]=16'h1030;
      mem[16'h050f]=16'h9220;
      mem[16'h0510]=16'h0654;
      mem[16'h0511]=16'hd552;
      mem[16'h0512]=16'h0841;
      mem[16'h0513]=16'h0831;
      mem[16'h0514]=16'h0170;
      mem[16'h0515]=16'hffbc;
      mem[16'h0516]=16'h01f0;
      mem[16'h0517]=16'h0002;
      mem[16'h0518]=16'h0002;
      mem[16'h0519]=16'h0002;
      mem[16'h051a]=16'h0a0d;
      mem[16'h051b]=16'h6e55;
      mem[16'h051c]=16'h7669;
      mem[16'h051d]=16'h7265;
      mem[16'h051e]=16'h6173;
      mem[16'h051f]=16'h206c;
      mem[16'h0520]=16'h6f4d;
      mem[16'h0521]=16'h696e;
      mem[16'h0522]=16'h6f74;
      mem[16'h0523]=16'h2072;
      mem[16'h0524]=16'h3848;
      mem[16'h0525]=16'h0d30;
      mem[16'h0526]=16'h000a;
      mem[16'h0527]=16'h205d;
      mem[16'h0528]=16'h4500;
      mem[16'h0529]=16'h7272;
      mem[16'h052a]=16'h726f;
      mem[16'h052b]=16'h6920;
      mem[16'h052c]=16'h6568;
      mem[16'h052d]=16'h0d78;
      mem[16'h052e]=16'h000a;
      mem[16'h052f]=16'h7245;
      mem[16'h0530]=16'h6f72;
      mem[16'h0531]=16'h2072;
      mem[16'h0532]=16'h7273;
      mem[16'h0533]=16'h6365;
      mem[16'h0534]=16'h0a0d;
      mem[16'h0535]=16'h4500;
      mem[16'h0536]=16'h7272;
      mem[16'h0537]=16'h726f;
      mem[16'h0538]=16'h0a0d;
      mem[16'h0539]=16'h2000;
      mem[16'h053a]=16'h003a;
      mem[16'h053b]=16'h3a20;
      mem[16'h053c]=16'h0020;
      mem[16'h053d]=16'h303a;
      mem[16'h053e]=16'h3030;
      mem[16'h053f]=16'h3030;
      mem[16'h0540]=16'h3030;
      mem[16'h0541]=16'h4631;
      mem[16'h0542]=16'h0d46;
      mem[16'h0543]=16'h000a;
      mem[16'h0544]=16'h3953;
      mem[16'h0545]=16'h3330;
      mem[16'h0546]=16'h3030;
      mem[16'h0547]=16'h3030;
      mem[16'h0548]=16'h4346;
      mem[16'h0549]=16'h0a0d;
      mem[16'h054a]=16'h4800;
      mem[16'h054b]=16'h3038;
      mem[16'h054c]=16'h3128;
      mem[16'h054d]=16'h2936;
      mem[16'h054e]=16'h0a0d;
      mem[16'h054f]=16'h4800;
      mem[16'h0550]=16'h3038;
      mem[16'h0551]=16'h3328;
      mem[16'h0552]=16'h2932;
      mem[16'h0553]=16'h0a0d;
      mem[16'h0554]=16'h5200;
      mem[16'h0555]=16'h5453;
      mem[16'h0556]=16'h3320;
      mem[16'h0557]=16'h4838;
      mem[16'h0558]=16'h0a0d;
      mem[16'h0559]=16'hff00;
      mem[16'h055a]=16'h0002;
      mem[16'h055b]=16'h0160;
      mem[16'h055c]=16'h0ac8;
      mem[16'h055d]=16'h01c0;
      mem[16'h055e]=16'h0170;
      mem[16'h055f]=16'hfff6;
      mem[16'h0560]=16'h03c0;
      mem[16'h0561]=16'h1000;
      mem[16'h0562]=16'h3b20;
      mem[16'h0563]=16'h0002;
      mem[16'h0564]=16'he222;
      mem[16'h0565]=16'h1001;
      mem[16'h0566]=16'h3b20;
      mem[16'h0567]=16'hd222;
      mem[16'h0568]=16'h0002;
      mem[16'h0569]=16'h1000;
      mem[16'h056a]=16'h3920;
      mem[16'h056b]=16'h0002;
      mem[16'h056c]=16'hffff;
      mem[16'h056d]=16'hffff;
      mem[16'h056e]=16'hffff;
      mem[16'h056f]=16'hffff;
      mem[16'h0570]=16'hffff;
      mem[16'h0571]=16'hffff;
      mem[16'h0572]=16'hffff;
      mem[16'h0573]=16'hffff;
      mem[16'h0574]=16'hffff;
      mem[16'h0575]=16'hffff;
      mem[16'h0576]=16'hffff;
      mem[16'h0577]=16'hffff;
      mem[16'h0578]=16'hffff;
      mem[16'h0579]=16'hffff;
      mem[16'h057a]=16'hffff;
      mem[16'h057b]=16'hffff;
      mem[16'h057c]=16'hffff;
      mem[16'h057d]=16'hffff;
      mem[16'h057e]=16'hffff;
      mem[16'h057f]=16'hffff;
      mem[16'h0580]=16'hffff;
      mem[16'h0581]=16'hffff;
      mem[16'h0582]=16'hffff;
      mem[16'h0583]=16'hffff;
      mem[16'h0584]=16'hffff;
      mem[16'h0585]=16'hffff;
      mem[16'h0586]=16'hffff;
      mem[16'h0587]=16'hffff;
      mem[16'h0588]=16'hffff;
      mem[16'h0589]=16'hffff;
      mem[16'h058a]=16'hffff;
      mem[16'h058b]=16'hffff;
      mem[16'h058c]=16'hffff;
      mem[16'h058d]=16'hffff;
      mem[16'h058e]=16'hffff;
      mem[16'h058f]=16'hffff;
      mem[16'h0590]=16'hffff;
      mem[16'h0591]=16'hffff;
      mem[16'h0592]=16'hffff;
      mem[16'h0593]=16'hffff;
      mem[16'h0594]=16'hffff;
      mem[16'h0595]=16'hffff;
      mem[16'h0596]=16'hffff;
      mem[16'h0597]=16'hffff;
      mem[16'h0598]=16'hffff;
      mem[16'h0599]=16'hffff;
      mem[16'h059a]=16'hffff;
      mem[16'h059b]=16'hffff;
      mem[16'h059c]=16'hffff;
      mem[16'h059d]=16'hffff;
      mem[16'h059e]=16'hffff;
      mem[16'h059f]=16'hffff;
      mem[16'h05a0]=16'hffff;
      mem[16'h05a1]=16'hffff;
      mem[16'h05a2]=16'hffff;
      mem[16'h05a3]=16'hffff;
      mem[16'h05a4]=16'hffff;
      mem[16'h05a5]=16'hffff;
      mem[16'h05a6]=16'hffff;
      mem[16'h05a7]=16'hffff;
      mem[16'h05a8]=16'hffff;
      mem[16'h05a9]=16'hffff;
      mem[16'h05aa]=16'hffff;
      mem[16'h05ab]=16'hffff;
      mem[16'h05ac]=16'hffff;
      mem[16'h05ad]=16'hffff;
      mem[16'h05ae]=16'hffff;
      mem[16'h05af]=16'hffff;
      mem[16'h05b0]=16'hffff;
      mem[16'h05b1]=16'hffff;
      mem[16'h05b2]=16'hffff;
      mem[16'h05b3]=16'hffff;
      mem[16'h05b4]=16'hffff;
      mem[16'h05b5]=16'hffff;
      mem[16'h05b6]=16'hffff;
      mem[16'h05b7]=16'hffff;
      mem[16'h05b8]=16'hffff;
      mem[16'h05b9]=16'hffff;
      mem[16'h05ba]=16'hffff;
      mem[16'h05bb]=16'hffff;
      mem[16'h05bc]=16'hffff;
      mem[16'h05bd]=16'hffff;
      mem[16'h05be]=16'hffff;
      mem[16'h05bf]=16'hffff;
      mem[16'h05c0]=16'hffff;
      mem[16'h05c1]=16'hffff;
      mem[16'h05c2]=16'hffff;
      mem[16'h05c3]=16'hffff;
      mem[16'h05c4]=16'hffff;
      mem[16'h05c5]=16'hffff;
      mem[16'h05c6]=16'hffff;
      mem[16'h05c7]=16'hffff;
      mem[16'h05c8]=16'hffff;
      mem[16'h05c9]=16'hffff;
      mem[16'h05ca]=16'hffff;
      mem[16'h05cb]=16'hffff;
      mem[16'h05cc]=16'hffff;
      mem[16'h05cd]=16'hffff;
      mem[16'h05ce]=16'hffff;
      mem[16'h05cf]=16'hffff;
      mem[16'h05d0]=16'hffff;
      mem[16'h05d1]=16'hffff;
      mem[16'h05d2]=16'hffff;
      mem[16'h05d3]=16'hffff;
      mem[16'h05d4]=16'hffff;
      mem[16'h05d5]=16'hffff;
      mem[16'h05d6]=16'hffff;
      mem[16'h05d7]=16'hffff;
      mem[16'h05d8]=16'hffff;
      mem[16'h05d9]=16'hffff;
      mem[16'h05da]=16'hffff;
      mem[16'h05db]=16'hffff;
      mem[16'h05dc]=16'hffff;
      mem[16'h05dd]=16'hffff;
      mem[16'h05de]=16'hffff;
      mem[16'h05df]=16'hffff;
      mem[16'h05e0]=16'hffff;
      mem[16'h05e1]=16'hffff;
      mem[16'h05e2]=16'hffff;
      mem[16'h05e3]=16'hffff;
      mem[16'h05e4]=16'hffff;
      mem[16'h05e5]=16'hffff;
      mem[16'h05e6]=16'hffff;
      mem[16'h05e7]=16'hffff;
      mem[16'h05e8]=16'hffff;
      mem[16'h05e9]=16'hffff;
      mem[16'h05ea]=16'hffff;
      mem[16'h05eb]=16'hffff;
      mem[16'h05ec]=16'hffff;
      mem[16'h05ed]=16'hffff;
      mem[16'h05ee]=16'hffff;
      mem[16'h05ef]=16'hffff;
      mem[16'h05f0]=16'hffff;
      mem[16'h05f1]=16'hffff;
      mem[16'h05f2]=16'hffff;
      mem[16'h05f3]=16'hffff;
      mem[16'h05f4]=16'hffff;
      mem[16'h05f5]=16'hffff;
      mem[16'h05f6]=16'hffff;
      mem[16'h05f7]=16'hffff;
      mem[16'h05f8]=16'hffff;
      mem[16'h05f9]=16'hffff;
      mem[16'h05fa]=16'hffff;
      mem[16'h05fb]=16'hffff;
      mem[16'h05fc]=16'hffff;
      mem[16'h05fd]=16'hffff;
      mem[16'h05fe]=16'hffff;
      mem[16'h05ff]=16'hffff;
      mem[16'h0600]=16'hffff;
      mem[16'h0601]=16'hffff;
      mem[16'h0602]=16'hffff;
      mem[16'h0603]=16'hffff;
      mem[16'h0604]=16'hffff;
      mem[16'h0605]=16'hffff;
      mem[16'h0606]=16'hffff;
      mem[16'h0607]=16'hffff;
      mem[16'h0608]=16'hffff;
      mem[16'h0609]=16'hffff;
      mem[16'h060a]=16'hffff;
      mem[16'h060b]=16'hffff;
      mem[16'h060c]=16'hffff;
      mem[16'h060d]=16'hffff;
      mem[16'h060e]=16'hffff;
      mem[16'h060f]=16'hffff;
      mem[16'h0610]=16'hffff;
      mem[16'h0611]=16'hffff;
      mem[16'h0612]=16'hffff;
      mem[16'h0613]=16'hffff;
      mem[16'h0614]=16'hffff;
      mem[16'h0615]=16'hffff;
      mem[16'h0616]=16'hffff;
      mem[16'h0617]=16'hffff;
      mem[16'h0618]=16'hffff;
      mem[16'h0619]=16'hffff;
      mem[16'h061a]=16'hffff;
      mem[16'h061b]=16'hffff;
      mem[16'h061c]=16'hffff;
      mem[16'h061d]=16'hffff;
      mem[16'h061e]=16'hffff;
      mem[16'h061f]=16'hffff;
      mem[16'h0620]=16'hffff;
      mem[16'h0621]=16'hffff;
      mem[16'h0622]=16'hffff;
      mem[16'h0623]=16'hffff;
      mem[16'h0624]=16'hffff;
      mem[16'h0625]=16'hffff;
      mem[16'h0626]=16'hffff;
      mem[16'h0627]=16'hffff;
      mem[16'h0628]=16'hffff;
      mem[16'h0629]=16'hffff;
      mem[16'h062a]=16'hffff;
      mem[16'h062b]=16'hffff;
      mem[16'h062c]=16'hffff;
      mem[16'h062d]=16'hffff;
      mem[16'h062e]=16'hffff;
      mem[16'h062f]=16'hffff;
      mem[16'h0630]=16'hffff;
      mem[16'h0631]=16'hffff;
      mem[16'h0632]=16'hffff;
      mem[16'h0633]=16'hffff;
      mem[16'h0634]=16'hffff;
      mem[16'h0635]=16'hffff;
      mem[16'h0636]=16'hffff;
      mem[16'h0637]=16'hffff;
      mem[16'h0638]=16'hffff;
      mem[16'h0639]=16'hffff;
      mem[16'h063a]=16'hffff;
      mem[16'h063b]=16'hffff;
      mem[16'h063c]=16'hffff;
      mem[16'h063d]=16'hffff;
      mem[16'h063e]=16'hffff;
      mem[16'h063f]=16'hffff;
      mem[16'h0640]=16'hffff;
      mem[16'h0641]=16'hffff;
      mem[16'h0642]=16'hffff;
      mem[16'h0643]=16'hffff;
      mem[16'h0644]=16'hffff;
      mem[16'h0645]=16'hffff;
      mem[16'h0646]=16'hffff;
      mem[16'h0647]=16'hffff;
      mem[16'h0648]=16'hffff;
      mem[16'h0649]=16'hffff;
      mem[16'h064a]=16'hffff;
      mem[16'h064b]=16'hffff;
      mem[16'h064c]=16'hffff;
      mem[16'h064d]=16'hffff;
      mem[16'h064e]=16'hffff;
      mem[16'h064f]=16'hffff;
      mem[16'h0650]=16'hffff;
      mem[16'h0651]=16'hffff;
      mem[16'h0652]=16'hffff;
      mem[16'h0653]=16'hffff;
      mem[16'h0654]=16'hffff;
      mem[16'h0655]=16'hffff;
      mem[16'h0656]=16'hffff;
      mem[16'h0657]=16'hffff;
      mem[16'h0658]=16'hffff;
      mem[16'h0659]=16'hffff;
      mem[16'h065a]=16'hffff;
      mem[16'h065b]=16'hffff;
      mem[16'h065c]=16'hffff;
      mem[16'h065d]=16'hffff;
      mem[16'h065e]=16'hffff;
      mem[16'h065f]=16'hffff;
      mem[16'h0660]=16'hffff;
      mem[16'h0661]=16'hffff;
      mem[16'h0662]=16'hffff;
      mem[16'h0663]=16'hffff;
      mem[16'h0664]=16'hffff;
      mem[16'h0665]=16'hffff;
      mem[16'h0666]=16'hffff;
      mem[16'h0667]=16'hffff;
      mem[16'h0668]=16'hffff;
      mem[16'h0669]=16'hffff;
      mem[16'h066a]=16'hffff;
      mem[16'h066b]=16'hffff;
      mem[16'h066c]=16'hffff;
      mem[16'h066d]=16'hffff;
      mem[16'h066e]=16'hffff;
      mem[16'h066f]=16'hffff;
      mem[16'h0670]=16'hffff;
      mem[16'h0671]=16'hffff;
      mem[16'h0672]=16'hffff;
      mem[16'h0673]=16'hffff;
      mem[16'h0674]=16'hffff;
      mem[16'h0675]=16'hffff;
      mem[16'h0676]=16'hffff;
      mem[16'h0677]=16'hffff;
      mem[16'h0678]=16'hffff;
      mem[16'h0679]=16'hffff;
      mem[16'h067a]=16'hffff;
      mem[16'h067b]=16'hffff;
      mem[16'h067c]=16'hffff;
      mem[16'h067d]=16'hffff;
      mem[16'h067e]=16'hffff;
      mem[16'h067f]=16'hffff;
      mem[16'h0680]=16'hffff;
      mem[16'h0681]=16'hffff;
      mem[16'h0682]=16'hffff;
      mem[16'h0683]=16'hffff;
      mem[16'h0684]=16'hffff;
      mem[16'h0685]=16'hffff;
      mem[16'h0686]=16'hffff;
      mem[16'h0687]=16'hffff;
      mem[16'h0688]=16'hffff;
      mem[16'h0689]=16'hffff;
      mem[16'h068a]=16'hffff;
      mem[16'h068b]=16'hffff;
      mem[16'h068c]=16'hffff;
      mem[16'h068d]=16'hffff;
      mem[16'h068e]=16'hffff;
      mem[16'h068f]=16'hffff;
      mem[16'h0690]=16'hffff;
      mem[16'h0691]=16'hffff;
      mem[16'h0692]=16'hffff;
      mem[16'h0693]=16'hffff;
      mem[16'h0694]=16'hffff;
      mem[16'h0695]=16'hffff;
      mem[16'h0696]=16'hffff;
      mem[16'h0697]=16'hffff;
      mem[16'h0698]=16'hffff;
      mem[16'h0699]=16'hffff;
      mem[16'h069a]=16'hffff;
      mem[16'h069b]=16'hffff;
      mem[16'h069c]=16'hffff;
      mem[16'h069d]=16'hffff;
      mem[16'h069e]=16'hffff;
      mem[16'h069f]=16'hffff;
      mem[16'h06a0]=16'hffff;
      mem[16'h06a1]=16'hffff;
      mem[16'h06a2]=16'hffff;
      mem[16'h06a3]=16'hffff;
      mem[16'h06a4]=16'hffff;
      mem[16'h06a5]=16'hffff;
      mem[16'h06a6]=16'hffff;
      mem[16'h06a7]=16'hffff;
      mem[16'h06a8]=16'hffff;
      mem[16'h06a9]=16'hffff;
      mem[16'h06aa]=16'hffff;
      mem[16'h06ab]=16'hffff;
      mem[16'h06ac]=16'hffff;
      mem[16'h06ad]=16'hffff;
      mem[16'h06ae]=16'hffff;
      mem[16'h06af]=16'hffff;
      mem[16'h06b0]=16'hffff;
      mem[16'h06b1]=16'hffff;
      mem[16'h06b2]=16'hffff;
      mem[16'h06b3]=16'hffff;
      mem[16'h06b4]=16'hffff;
      mem[16'h06b5]=16'hffff;
      mem[16'h06b6]=16'hffff;
      mem[16'h06b7]=16'hffff;
      mem[16'h06b8]=16'hffff;
      mem[16'h06b9]=16'hffff;
      mem[16'h06ba]=16'hffff;
      mem[16'h06bb]=16'hffff;
      mem[16'h06bc]=16'hffff;
      mem[16'h06bd]=16'hffff;
      mem[16'h06be]=16'hffff;
      mem[16'h06bf]=16'hffff;
      mem[16'h06c0]=16'hffff;
      mem[16'h06c1]=16'hffff;
      mem[16'h06c2]=16'hffff;
      mem[16'h06c3]=16'hffff;
      mem[16'h06c4]=16'hffff;
      mem[16'h06c5]=16'hffff;
      mem[16'h06c6]=16'hffff;
      mem[16'h06c7]=16'hffff;
      mem[16'h06c8]=16'hffff;
      mem[16'h06c9]=16'hffff;
      mem[16'h06ca]=16'hffff;
      mem[16'h06cb]=16'hffff;
      mem[16'h06cc]=16'hffff;
      mem[16'h06cd]=16'hffff;
      mem[16'h06ce]=16'hffff;
      mem[16'h06cf]=16'hffff;
      mem[16'h06d0]=16'hffff;
      mem[16'h06d1]=16'hffff;
      mem[16'h06d2]=16'hffff;
      mem[16'h06d3]=16'hffff;
      mem[16'h06d4]=16'hffff;
      mem[16'h06d5]=16'hffff;
      mem[16'h06d6]=16'hffff;
      mem[16'h06d7]=16'hffff;
      mem[16'h06d8]=16'hffff;
      mem[16'h06d9]=16'hffff;
      mem[16'h06da]=16'hffff;
      mem[16'h06db]=16'hffff;
      mem[16'h06dc]=16'hffff;
      mem[16'h06dd]=16'hffff;
      mem[16'h06de]=16'hffff;
      mem[16'h06df]=16'hffff;
      mem[16'h06e0]=16'hffff;
      mem[16'h06e1]=16'hffff;
      mem[16'h06e2]=16'hffff;
      mem[16'h06e3]=16'hffff;
      mem[16'h06e4]=16'hffff;
      mem[16'h06e5]=16'hffff;
      mem[16'h06e6]=16'hffff;
      mem[16'h06e7]=16'hffff;
      mem[16'h06e8]=16'hffff;
      mem[16'h06e9]=16'hffff;
      mem[16'h06ea]=16'hffff;
      mem[16'h06eb]=16'hffff;
      mem[16'h06ec]=16'hffff;
      mem[16'h06ed]=16'hffff;
      mem[16'h06ee]=16'hffff;
      mem[16'h06ef]=16'hffff;
      mem[16'h06f0]=16'hffff;
      mem[16'h06f1]=16'hffff;
      mem[16'h06f2]=16'hffff;
      mem[16'h06f3]=16'hffff;
      mem[16'h06f4]=16'hffff;
      mem[16'h06f5]=16'hffff;
      mem[16'h06f6]=16'hffff;
      mem[16'h06f7]=16'hffff;
      mem[16'h06f8]=16'hffff;
      mem[16'h06f9]=16'hffff;
      mem[16'h06fa]=16'hffff;
      mem[16'h06fb]=16'hffff;
      mem[16'h06fc]=16'hffff;
      mem[16'h06fd]=16'hffff;
      mem[16'h06fe]=16'hffff;
      mem[16'h06ff]=16'hffff;
      mem[16'h0700]=16'hffff;
      mem[16'h0701]=16'hffff;
      mem[16'h0702]=16'hffff;
      mem[16'h0703]=16'hffff;
      mem[16'h0704]=16'hffff;
      mem[16'h0705]=16'hffff;
      mem[16'h0706]=16'hffff;
      mem[16'h0707]=16'hffff;
      mem[16'h0708]=16'hffff;
      mem[16'h0709]=16'hffff;
      mem[16'h070a]=16'hffff;
      mem[16'h070b]=16'hffff;
      mem[16'h070c]=16'hffff;
      mem[16'h070d]=16'hffff;
      mem[16'h070e]=16'hffff;
      mem[16'h070f]=16'hffff;
      mem[16'h0710]=16'hffff;
      mem[16'h0711]=16'hffff;
      mem[16'h0712]=16'hffff;
      mem[16'h0713]=16'hffff;
      mem[16'h0714]=16'hffff;
      mem[16'h0715]=16'hffff;
      mem[16'h0716]=16'hffff;
      mem[16'h0717]=16'hffff;
      mem[16'h0718]=16'hffff;
      mem[16'h0719]=16'hffff;
      mem[16'h071a]=16'hffff;
      mem[16'h071b]=16'hffff;
      mem[16'h071c]=16'hffff;
      mem[16'h071d]=16'hffff;
      mem[16'h071e]=16'hffff;
      mem[16'h071f]=16'hffff;
      mem[16'h0720]=16'hffff;
      mem[16'h0721]=16'hffff;
      mem[16'h0722]=16'hffff;
      mem[16'h0723]=16'hffff;
      mem[16'h0724]=16'hffff;
      mem[16'h0725]=16'hffff;
      mem[16'h0726]=16'hffff;
      mem[16'h0727]=16'hffff;
      mem[16'h0728]=16'hffff;
      mem[16'h0729]=16'hffff;
      mem[16'h072a]=16'hffff;
      mem[16'h072b]=16'hffff;
      mem[16'h072c]=16'hffff;
      mem[16'h072d]=16'hffff;
      mem[16'h072e]=16'hffff;
      mem[16'h072f]=16'hffff;
      mem[16'h0730]=16'hffff;
      mem[16'h0731]=16'hffff;
      mem[16'h0732]=16'hffff;
      mem[16'h0733]=16'hffff;
      mem[16'h0734]=16'hffff;
      mem[16'h0735]=16'hffff;
      mem[16'h0736]=16'hffff;
      mem[16'h0737]=16'hffff;
      mem[16'h0738]=16'hffff;
      mem[16'h0739]=16'hffff;
      mem[16'h073a]=16'hffff;
      mem[16'h073b]=16'hffff;
      mem[16'h073c]=16'hffff;
      mem[16'h073d]=16'hffff;
      mem[16'h073e]=16'hffff;
      mem[16'h073f]=16'hffff;
      mem[16'h0740]=16'hffff;
      mem[16'h0741]=16'hffff;
      mem[16'h0742]=16'hffff;
      mem[16'h0743]=16'hffff;
      mem[16'h0744]=16'hffff;
      mem[16'h0745]=16'hffff;
      mem[16'h0746]=16'hffff;
      mem[16'h0747]=16'hffff;
      mem[16'h0748]=16'hffff;
      mem[16'h0749]=16'hffff;
      mem[16'h074a]=16'hffff;
      mem[16'h074b]=16'hffff;
      mem[16'h074c]=16'hffff;
      mem[16'h074d]=16'hffff;
      mem[16'h074e]=16'hffff;
      mem[16'h074f]=16'hffff;
      mem[16'h0750]=16'hffff;
      mem[16'h0751]=16'hffff;
      mem[16'h0752]=16'hffff;
      mem[16'h0753]=16'hffff;
      mem[16'h0754]=16'hffff;
      mem[16'h0755]=16'hffff;
      mem[16'h0756]=16'hffff;
      mem[16'h0757]=16'hffff;
      mem[16'h0758]=16'hffff;
      mem[16'h0759]=16'hffff;
      mem[16'h075a]=16'hffff;
      mem[16'h075b]=16'hffff;
      mem[16'h075c]=16'hffff;
      mem[16'h075d]=16'hffff;
      mem[16'h075e]=16'hffff;
      mem[16'h075f]=16'hffff;
      mem[16'h0760]=16'hffff;
      mem[16'h0761]=16'hffff;
      mem[16'h0762]=16'hffff;
      mem[16'h0763]=16'hffff;
      mem[16'h0764]=16'hffff;
      mem[16'h0765]=16'hffff;
      mem[16'h0766]=16'hffff;
      mem[16'h0767]=16'hffff;
      mem[16'h0768]=16'hffff;
      mem[16'h0769]=16'hffff;
      mem[16'h076a]=16'hffff;
      mem[16'h076b]=16'hffff;
      mem[16'h076c]=16'hffff;
      mem[16'h076d]=16'hffff;
      mem[16'h076e]=16'hffff;
      mem[16'h076f]=16'hffff;
      mem[16'h0770]=16'hffff;
      mem[16'h0771]=16'hffff;
      mem[16'h0772]=16'hffff;
      mem[16'h0773]=16'hffff;
      mem[16'h0774]=16'hffff;
      mem[16'h0775]=16'hffff;
      mem[16'h0776]=16'hffff;
      mem[16'h0777]=16'hffff;
      mem[16'h0778]=16'hffff;
      mem[16'h0779]=16'hffff;
      mem[16'h077a]=16'hffff;
      mem[16'h077b]=16'hffff;
      mem[16'h077c]=16'hffff;
      mem[16'h077d]=16'hffff;
      mem[16'h077e]=16'hffff;
      mem[16'h077f]=16'hffff;
      mem[16'h0780]=16'hffff;
      mem[16'h0781]=16'hffff;
      mem[16'h0782]=16'hffff;
      mem[16'h0783]=16'hffff;
      mem[16'h0784]=16'hffff;
      mem[16'h0785]=16'hffff;
      mem[16'h0786]=16'hffff;
      mem[16'h0787]=16'hffff;
      mem[16'h0788]=16'hffff;
      mem[16'h0789]=16'hffff;
      mem[16'h078a]=16'hffff;
      mem[16'h078b]=16'hffff;
      mem[16'h078c]=16'hffff;
      mem[16'h078d]=16'hffff;
      mem[16'h078e]=16'hffff;
      mem[16'h078f]=16'hffff;
      mem[16'h0790]=16'hffff;
      mem[16'h0791]=16'hffff;
      mem[16'h0792]=16'hffff;
      mem[16'h0793]=16'hffff;
      mem[16'h0794]=16'hffff;
      mem[16'h0795]=16'hffff;
      mem[16'h0796]=16'hffff;
      mem[16'h0797]=16'hffff;
      mem[16'h0798]=16'hffff;
      mem[16'h0799]=16'hffff;
      mem[16'h079a]=16'hffff;
      mem[16'h079b]=16'hffff;
      mem[16'h079c]=16'hffff;
      mem[16'h079d]=16'hffff;
      mem[16'h079e]=16'hffff;
      mem[16'h079f]=16'hffff;
      mem[16'h07a0]=16'hffff;
      mem[16'h07a1]=16'hffff;
      mem[16'h07a2]=16'hffff;
      mem[16'h07a3]=16'hffff;
      mem[16'h07a4]=16'hffff;
      mem[16'h07a5]=16'hffff;
      mem[16'h07a6]=16'hffff;
      mem[16'h07a7]=16'hffff;
      mem[16'h07a8]=16'hffff;
      mem[16'h07a9]=16'hffff;
      mem[16'h07aa]=16'hffff;
      mem[16'h07ab]=16'hffff;
      mem[16'h07ac]=16'hffff;
      mem[16'h07ad]=16'hffff;
      mem[16'h07ae]=16'hffff;
      mem[16'h07af]=16'hffff;
      mem[16'h07b0]=16'hffff;
      mem[16'h07b1]=16'hffff;
      mem[16'h07b2]=16'hffff;
      mem[16'h07b3]=16'hffff;
      mem[16'h07b4]=16'hffff;
      mem[16'h07b5]=16'hffff;
      mem[16'h07b6]=16'hffff;
      mem[16'h07b7]=16'hffff;
      mem[16'h07b8]=16'hffff;
      mem[16'h07b9]=16'hffff;
      mem[16'h07ba]=16'hffff;
      mem[16'h07bb]=16'hffff;
      mem[16'h07bc]=16'hffff;
      mem[16'h07bd]=16'hffff;
      mem[16'h07be]=16'hffff;
      mem[16'h07bf]=16'hffff;
      mem[16'h07c0]=16'hffff;
      mem[16'h07c1]=16'hffff;
      mem[16'h07c2]=16'hffff;
      mem[16'h07c3]=16'hffff;
      mem[16'h07c4]=16'hffff;
      mem[16'h07c5]=16'hffff;
      mem[16'h07c6]=16'hffff;
      mem[16'h07c7]=16'hffff;
      mem[16'h07c8]=16'hffff;
      mem[16'h07c9]=16'hffff;
      mem[16'h07ca]=16'hffff;
      mem[16'h07cb]=16'hffff;
      mem[16'h07cc]=16'hffff;
      mem[16'h07cd]=16'hffff;
      mem[16'h07ce]=16'hffff;
      mem[16'h07cf]=16'hffff;
      mem[16'h07d0]=16'hffff;
      mem[16'h07d1]=16'hffff;
      mem[16'h07d2]=16'hffff;
      mem[16'h07d3]=16'hffff;
      mem[16'h07d4]=16'hffff;
      mem[16'h07d5]=16'hffff;
      mem[16'h07d6]=16'hffff;
      mem[16'h07d7]=16'hffff;
      mem[16'h07d8]=16'hffff;
      mem[16'h07d9]=16'hffff;
      mem[16'h07da]=16'hffff;
      mem[16'h07db]=16'hffff;
      mem[16'h07dc]=16'hffff;
      mem[16'h07dd]=16'hffff;
      mem[16'h07de]=16'hffff;
      mem[16'h07df]=16'hffff;
      mem[16'h07e0]=16'hffff;
      mem[16'h07e1]=16'hffff;
      mem[16'h07e2]=16'hffff;
      mem[16'h07e3]=16'hffff;
      mem[16'h07e4]=16'hffff;
      mem[16'h07e5]=16'hffff;
      mem[16'h07e6]=16'hffff;
      mem[16'h07e7]=16'hffff;
      mem[16'h07e8]=16'hffff;
      mem[16'h07e9]=16'hffff;
      mem[16'h07ea]=16'hffff;
      mem[16'h07eb]=16'hffff;
      mem[16'h07ec]=16'hffff;
      mem[16'h07ed]=16'hffff;
      mem[16'h07ee]=16'hffff;
      mem[16'h07ef]=16'hffff;
      mem[16'h07f0]=16'hffff;
      mem[16'h07f1]=16'hffff;
      mem[16'h07f2]=16'hffff;
      mem[16'h07f3]=16'hffff;
      mem[16'h07f4]=16'hffff;
      mem[16'h07f5]=16'hffff;
      mem[16'h07f6]=16'hffff;
      mem[16'h07f7]=16'hffff;
      mem[16'h07f8]=16'hffff;
      mem[16'h07f9]=16'hffff;
      mem[16'h07fa]=16'hffff;
      mem[16'h07fb]=16'hffff;
      mem[16'h07fc]=16'hffff;
      mem[16'h07fd]=16'hffff;
      mem[16'h07fe]=16'hffff;
      mem[16'h07ff]=16'hffff;
      mem[16'h0800]=16'h0000;
end
