      mem['h0800] = 'h0444;  // I_SRA_R_I(4, 4)
      mem['h0801] = 'h0455;  // I_SRA_R_I(5, FRACBITS - 4)
      mem['h0802] = 'ha245;  // I_MUL(2, 4, 5)
      mem['h0803] = 'h0002;  // I_RET()
      mem['h0804] = 'h0178;  // I_LD_RW_I(8)
      mem['h0805] = 'h000a;  // 10
      mem['h0806] = 'hf448;  // I_CP(4, 4, 8)
      mem['h0807] = 'h0178;  // I_LD_RW_I(8)
      mem['h0808] = 'h0004;  // 4
      mem['h0809] = 'h03d8;  // I_JR_C(8)
      mem['h080a] = 'h0847;  // I_ADD_R_I(4, 7)
      mem['h080b] = 'h0178;  // I_LD_RW_I(8)
      mem['h080c] = 'h0030;  // 48
      mem['h080d] = 'h8448;  // I_ADD(4, 4, 8)
      mem['h080e] = 'h0178;  // I_LD_RW_I(8)
      mem['h080f] = 'h0000;  // 'h0000
      mem['h0810] = 'h3948;  // I_OUTB(8, 4)
      mem['h0811] = 'h0002;  // I_RET()
      mem['h0000] = 'h0170;  // I_LD_RW_I(0)
      mem['h0001] = 'h0000;  // 'h0000
      mem['h0002] = 'h3f20;  // I_LD_R_R(reg_sp, 0)
      mem['h0003] = 'h017e;  // I_LD_RW_I(CA)
      mem['h0004] = 'hfc7f;  // CA0
      mem['h0005] = 'h017f;  // I_LD_RW_I(CB)
      mem['h0006] = 'hfe08;  // CB0
      mem['h0007] = 'h0177;  // I_LD_RW_I(Y)
      mem['h0008] = 'h0018;  // HEIGHT
      mem['h0009] = 'h0871;  // I_ADD_R_I(Y, 1)
      mem['h000a] = 'h017e;  // I_LD_RW_I(CA)
      mem['h000b] = 'hfc7f;  // CA0
      mem['h000c] = 'h0176;  // I_LD_RW_I(X)
      mem['h000d] = 'h004e;  // WIDTH
      mem['h000e] = 'h0861;  // I_ADD_R_I(X, 1)
      mem['h000f] = 'h3cec;  // I_LD_R_R(A, CA)
      mem['h0010] = 'h3cfd;  // I_LD_R_R(B, CB)
      mem['h0011] = 'hebbb;  // I_XOR(I, I, I)
      mem['h0012] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h0013] = 'h3cc5;  // I_LD_R_R(5, A)
      mem['h0014] = 'h0170;  // I_LD_RW_I(0)
      mem['h0015] = 'h1000;  // label_fp_mul
      mem['h0016] = 'h01c0;  // I_CALL_R(0)
      mem['h0017] = 'h3c23;  // I_LD_R_R(T, 2)
      mem['h0018] = 'h3cd4;  // I_LD_R_R(4, B)
      mem['h0019] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h001a] = 'h0170;  // I_LD_RW_I(0)
      mem['h001b] = 'h1000;  // label_fp_mul
      mem['h001c] = 'h01c0;  // I_CALL_R(0)
      mem['h001d] = 'h9332;  // I_SUB(T, T, 2)
      mem['h001e] = 'h833e;  // I_ADD(T, T, CA)
      mem['h001f] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h0020] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h0021] = 'h0170;  // I_LD_RW_I(0)
      mem['h0022] = 'h1000;  // label_fp_mul
      mem['h0023] = 'h01c0;  // I_CALL_R(0)
      mem['h0024] = 'h0621;  // I_SL_R_I(2, 1)
      mem['h0025] = 'h8d2f;  // I_ADD(B, 2, CB)
      mem['h0026] = 'h3c3c;  // I_LD_R_R(A, T)
      mem['h0027] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h0028] = 'h3cc5;  // I_LD_R_R(5, A)
      mem['h0029] = 'h0170;  // I_LD_RW_I(0)
      mem['h002a] = 'h1000;  // label_fp_mul
      mem['h002b] = 'h01c0;  // I_CALL_R(0)
      mem['h002c] = 'h3c23;  // I_LD_R_R(T, 2)
      mem['h002d] = 'h3cd4;  // I_LD_R_R(4, B)
      mem['h002e] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h002f] = 'h0170;  // I_LD_RW_I(0)
      mem['h0030] = 'h1000;  // label_fp_mul
      mem['h0031] = 'h01c0;  // I_CALL_R(0)
      mem['h0032] = 'h8332;  // I_ADD(T, T, 2)
      mem['h0033] = 'h0170;  // I_LD_RW_I(0)
      mem['h0034] = 'h0800;  // FP4_0
      mem['h0035] = 'hf303;  // I_CP(T, 0, T)
      mem['h0036] = 'h0170;  // I_LD_RW_I(0)
      mem['h0037] = 'h0010;  // 16
      mem['h0038] = 'h0390;  // I_JR_NC(0)
      mem['h0039] = 'h3cb4;  // I_LD_R_R(4, I)
      mem['h003a] = 'h0170;  // I_LD_RW_I(0)
      mem['h003b] = 'h1008;  // label_put_pixel
      mem['h003c] = 'h01c0;  // I_CALL_R(0)
      mem['h003d] = 'h0170;  // I_LD_RW_I(0)
      mem['h003f] = 'h01e0;  // I_JP_R(0)
      mem['h0040] = 'h08b1;  // I_ADD_R_I(I, 1)
      mem['h0041] = 'h0170;  // I_LD_RW_I(0)
      mem['h0042] = 'h0010;  // 16
      mem['h0043] = 'hfbb0;  // I_CP(I, I, 0)
      mem['h0044] = 'h0170;  // I_LD_RW_I(0)
      mem['h0045] = 'h0024;  // label_loop_i
      mem['h0046] = 'h0350;  // I_JP_C(0)
      mem['h0047] = 'h0171;  // I_LD_RW_I(1)
      mem['h0048] = 'h0000;  // 'h0000
      mem['h0049] = 'h1020;  // I_LD_RL_I(0, 'h20)
      mem['h004a] = 'h3901;  // I_OUTB(1, 0)
      mem['h003e] = 'h0096;  // addr
      mem['h004b] = 'h0170;  // I_LD_RW_I(0)
      mem['h004c] = 'h0017;  // FP0_0458
      mem['h004d] = 'h8ee0;  // I_ADD(CA, CA, 0)
      mem['h004e] = 'h0961;  // I_SUB_R_I(X, 1)
      mem['h004f] = 'h0170;  // I_LD_RW_I(0)
      mem['h0050] = 'h001e;  // label_loop_x
      mem['h0051] = 'h0300;  // I_JP_NZ(0)
      mem['h0052] = 'h0170;  // I_LD_RW_I(0)
      mem['h0053] = 'h002a;  // FP0_0833
      mem['h0054] = 'h8ff0;  // I_ADD(CB, CB, 0)
      mem['h0055] = 'h0171;  // I_LD_RW_I(1)
      mem['h0056] = 'h0000;  // 'h0000
      mem['h0057] = 'h100d;  // I_LD_RL_I(0, 'h0d)
      mem['h0058] = 'h3901;  // I_OUTB(1, 0)
      mem['h0059] = 'h100a;  // I_LD_RL_I(0, 'h0a)
      mem['h005a] = 'h3901;  // I_OUTB(1, 0)
      mem['h005b] = 'h0971;  // I_SUB_R_I(Y, 1)
      mem['h005c] = 'h0170;  // I_LD_RW_I(0)
      mem['h005d] = 'h0014;  // label_loop_y
      mem['h005e] = 'h0300;  // I_JP_NZ(0)
      mem['h005f] = 'h0001;  // I_HALT()
