   `include "h80cpu.svh"
   `include "h80cpu_instmacros.svh"
   initial begin
      mem['h0800] = 'h0444;  // I_SRA_R_I(4, 4)
      mem['h0801] = 'h0455;  // I_SRA_R_I(5, FRACBITS - 4)
      mem['h0802] = 'ha245;  // I_MUL(2, 4, 5)
      mem['h0803] = 'h0002;  // I_RET()
      mem['h0804] = 'h0168;  // I_LD_RW_I(8)
      mem['h0805] = 'h000a;  // 10
      mem['h0806] = 'hf448;  // I_CP(4, 4, 8)
      mem['h0807] = 'h0168;  // I_LD_RW_I(8)
      mem['h0808] = 'h0004;  // 4
      mem['h0809] = 'h03d8;  // I_JR_C(8)
      mem['h080a] = 'h0847;  // I_ADD_R_I(4, 7)
      mem['h080b] = 'h0168;  // I_LD_RW_I(8)
      mem['h080c] = 'h0030;  // 48
      mem['h080d] = 'h8448;  // I_ADD(4, 4, 8)
      mem['h080e] = 'h0168;  // I_LD_RW_I(8)
      mem['h080f] = 'h0000;
      mem['h0810] = 'h3948;  // I_OUTB(8, 4)
      mem['h0811] = 'h0002;  // I_RET()
      mem['h0000] = 'h0160;  // I_LD_RW_I(0)
      mem['h0001] = 'h4000;  // 'h4000
      mem['h0002] = 'h3f20;  // I_LD_R_R(reg_sp, 0)
      mem['h0003] = 'h017f;  // I_LD_RW_SI(CB)
      mem['h0004] = 'hfe08;  // CB0
      mem['h0005] = 'h0177;  // I_LD_RW_SI(Y)
      mem['h0006] = 'h0018;
      mem['h0007] = 'h0871;
      mem['h0008] = 'h017e;  // I_LD_RW_SI(CA)
      mem['h0009] = 'hfc7f;  // CA0
      mem['h000a] = 'h0176;  // I_LD_RW_SI(X)
      mem['h000b] = 'h004e;
      mem['h000c] = 'h0861;  // I_ADD_R_I(X, 1)
      mem['h000d] = 'h3cec;  // I_LD_R_R(A, CA)
      mem['h000e] = 'h3cfd;  // I_LD_R_R(B, CB)
      mem['h000f] = 'hebbb;  // I_XOR(I, I, I)
      mem['h0010] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h0011] = 'h3cc5;  // I_LD_R_R(5, A)
      mem['h0012] = 'h0160;  // I_LD_RW_I(0)
      mem['h0013] = 'h1000;
      mem['h0014] = 'h01c0;  // I_CALL_R(0)
      mem['h0015] = 'h3c23;  // I_LD_R_R(T, 2)
      mem['h0016] = 'h3cd4;  // I_LD_R_R(4, B)
      mem['h0017] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h0018] = 'h0160;  // I_LD_RW_I(0)
      mem['h0019] = 'h1000;
      mem['h001a] = 'h01c0;  // I_CALL_R(0)
      mem['h001b] = 'h9332;  // I_SUB(T, T, 2)
      mem['h001c] = 'h833e;  // I_ADD(T, T, CA)
      mem['h001d] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h001e] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h001f] = 'h0160;  // I_LD_RW_I(0)
      mem['h0020] = 'h1000;
      mem['h0021] = 'h01c0;  // I_CALL_R(0)
      mem['h0022] = 'h0621;  // I_SL_R_I(2, 1)
      mem['h0023] = 'h8d2f;  // I_ADD(B, 2, CB)
      mem['h0024] = 'h3c3c;  // I_LD_R_R(A, T)
      mem['h0025] = 'h3cc4;  // I_LD_R_R(4, A)
      mem['h0026] = 'h3cc5;  // I_LD_R_R(5, A)
      mem['h0027] = 'h0160;  // I_LD_RW_I(0)
      mem['h0028] = 'h1000;
      mem['h0029] = 'h01c0;  // I_CALL_R(0)
      mem['h002a] = 'h3c23;  // I_LD_R_R(T, 2)
      mem['h002b] = 'h3cd4;  // I_LD_R_R(4, B)
      mem['h002c] = 'h3cd5;  // I_LD_R_R(5, B)
      mem['h002d] = 'h0160;  // I_LD_RW_I(0)
      mem['h002e] = 'h1000;
      mem['h002f] = 'h01c0;  // I_CALL_R(0)
      mem['h0030] = 'h8332;  // I_ADD(T, T, 2)
      mem['h0031] = 'h0160;  // I_LD_RW_I(0)
      mem['h0032] = 'h0800;
      mem['h0033] = 'h0161;  // I_LD_RW_I(1)
      mem['h0034] = 'h0010;
      mem['h0035] = 'hf303;  // I_CP(T, 0, T)
      mem['h0036] = 'h0391;  // I_JR_NC(1)
      mem['h0037] = 'h3cb4;  // I_LD_R_R(4, I)
      mem['h0038] = 'h0160;  // I_LD_RW_I(0)
      mem['h0039] = 'h1008;
      mem['h003a] = 'h01c0;  // I_CALL_R(0)
      mem['h003b] = 'h0160;  // I_LD_RW_I(0)
      mem['h003c] = 'h0092;
      mem['h003d] = 'h01e0;  // I_JP_R(0)
      mem['h003e] = 'h08b1;  // I_ADD_R_I(I, 1)
      mem['h003f] = 'h0160;  // I_LD_RW_I(0)
      mem['h0040] = 'h0010;
      mem['h0041] = 'h0161;  // I_LD_RW_I(1)
      mem['h0042] = 'h0020;
      mem['h0043] = 'hfbb0;  // I_CP(I, I, 0)
      mem['h0044] = 'h0351;  // I_JP_C(1)
      mem['h0045] = 'h0161;  // I_LD_RW_I(1)
      mem['h0046] = 'h0000;
      mem['h0047] = 'h1020;  // I_LD_RB_I(0, 'h20)
      mem['h0048] = 'h3901;  // I_OUTB(1, 0)
      mem['h0049] = 'h0160;  // I_LD_RW_I(0)
      mem['h004a] = 'h0017;
      mem['h004b] = 'h8ee0;  // I_ADD(CA, CA, 0)
      mem['h004c] = 'h0160;  // I_LD_RW_I(0)
      mem['h004d] = 'h001a;
      mem['h004e] = 'h0961;  // I_SUB_R_I(X, 1)
      mem['h004f] = 'h0300;  // I_JP_NZ(0)
      mem['h0050] = 'h0170;  // I_LD_RW_SI(0)
      mem['h0051] = 'h002a;
      mem['h0052] = 'h8ff0;  // I_ADD(CB, CB, 0)
      mem['h0053] = 'h0161;  // I_LD_RW_I(1)
      mem['h0054] = 'h0000;
      mem['h0055] = 'h100d;  // I_LD_RB_I(0, 'h0d)
      mem['h0056] = 'h3901;  // I_OUTB(1, 0)
      mem['h0057] = 'h100a;  // I_LD_RB_I(0, 'h0a)
      mem['h0058] = 'h3901;  // I_OUTB(1, 0)
      mem['h0059] = 'h0160;  // I_LD_RW_I(0)
      mem['h005a] = 'h0010;
      mem['h005b] = 'h0971;  // I_SUB_R_I(Y, 1)
      mem['h005c] = 'h0300;  // I_JP_NZ(0)
      mem['h005d] = 'h0001;  // I_HALT()
   end
